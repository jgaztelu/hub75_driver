module bulbasaur_rom #(
    parameter hpixel_p = 64,
    parameter vpixel_p = 64,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p * vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
) (

    // Clock and reset
    input logic clk,
    input logic rst_n,

    /* Pixel read interface */
    input logic [addr_width_p-1:0] i_rd_addr,
    output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
);

  localparam bulbasaur_rom_buf[frame_size_p-1:0] = {
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454271,
    8454271,
    8454271,
    8454271,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454271,
    8454271,
    8454271,
    8454271,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454271,
    8454271,
    8454271,
    8454271,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454271,
    8454271,
    8454271,
    8454271,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8454269,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454271,
    8454271,
    8454271,
    8454271,
    8454269,
    8454269,
    8454271,
    8454271,
    8454271,
    8454271,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454273,
    8454271,
    8454271,
    8454271,
    8454271,
    8454269,
    8454269,
    8454271,
    8454271,
    8454271,
    8454271,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454271,
    8454271,
    8454271,
    8454271,
    8454273,
    8454273,
    8454271,
    8454271,
    8323199,
    8323199,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454271,
    8454271,
    8454271,
    8454271,
    8454273,
    8454273,
    8454271,
    8454271,
    8323199,
    8323199,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454271,
    8454271,
    8454271,
    8454271,
    8454271,
    8454271,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454271,
    8454271,
    8454271,
    8454271,
    8454271,
    8454271,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454269,
    8454269,
    8454269,
    8454269,
    8454271,
    8454271,
    8323199,
    8323199,
    8257663,
    8257663,
    8257663,
    8126847,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454269,
    8454269,
    8454269,
    8454269,
    8454271,
    8454271,
    8323199,
    8323199,
    8257663,
    8257663,
    8126847,
    8126847,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454269,
    8454269,
    8454269,
    8454269,
    8454271,
    8454271,
    8323199,
    8323199,
    8257663,
    8257663,
    8257663,
    8257663,
    8257665,
    8257665,
    8257665,
    8257665,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454269,
    8454269,
    8454269,
    8454269,
    8454271,
    8454271,
    8323199,
    8323199,
    8257663,
    8257663,
    8257663,
    8257663,
    8257665,
    8257665,
    8257665,
    8257665,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454269,
    8454269,
    8454269,
    8454269,
    8454271,
    8454271,
    8323199,
    8323199,
    8257663,
    8257663,
    8257663,
    8257663,
    8257665,
    8257665,
    8257665,
    8257665,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454269,
    8454269,
    8454269,
    8454269,
    8454271,
    8454271,
    8323199,
    8323199,
    8257663,
    8257663,
    8257663,
    8257663,
    8257665,
    8257665,
    8257665,
    8257665,
    8126847,
    8126847,
    8323199,
    8323199,
    8257663,
    8257663,
    8454271,
    8585343,
    8454273,
    8454273,
    8454271,
    8323197,
    8257917,
    8192125,
    8585603,
    8585345,
    8323201,
    8257663,
    8257663,
    8257917,
    8257917,
    8257915,
    8257915,
    8127097,
    7931253,
    8062071,
    8323195,
    8454271,
    8323201,
    8257665,
    8126847,
    8126847,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8126847,
    7799935,
    7930749,
    8585341,
    8585341,
    8127101,
    8127101,
    8650877,
    8847489,
    8781959,
    8650885,
    8585343,
    8323195,
    8522368,
    7798902,
    9044104,
    9109641,
    8980620,
    8389765,
    8192894,
    8061306,
    7864434,
    7995761,
    8390772,
    7603303,
    7542378,
    7080291,
    8192626,
    8257656,
    8257669,
    8061317,
    8061569,
    8126847,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8257663,
    7930751,
    8061567,
    8650879,
    8650879,
    8061567,
    8061567,
    8585343,
    8781955,
    8781959,
    8650887,
    8454273,
    8061051,
    7667828,
    7733365,
    8586115,
    7995517,
    7473530,
    6292074,
    6489449,
    7542389,
    6753123,
    7674477,
    7279973,
    6427990,
    5645644,
    6961250,
    6623838,
    6619233,
    7538042,
    7799935,
    8061821,
    8127101,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257665,
    8257665,
    8323201,
    8323201,
    8323201,
    8323201,
    8257665,
    8323201,
    8650883,
    8585347,
    8061315,
    7931012,
    8126597,
    8323205,
    8585349,
    8454277,
    8126599,
    8323719,
    8651910,
    8259198,
    6817133,
    6493549,
    5841513,
    4923741,
    4726870,
    4924245,
    4463944,
    5122126,
    4595780,
    5850966,
    4017977,
    9348237,
    985362,
    2687020,
    6295388,
    7604591,
    7931253,
    8127097,
    8257917,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257665,
    8257665,
    8323201,
    8323201,
    8323201,
    8323201,
    8257665,
    8323201,
    8323203,
    8323203,
    7864449,
    7996292,
    8061317,
    8126851,
    8323201,
    8323201,
    8061315,
    7734655,
    7670904,
    6557540,
    5382232,
    7889025,
    7631237,
    7962250,
    6909558,
    4738897,
    4870733,
    4673350,
    4739397,
    9414795,
    5342795,
    5409617,
    3824705,
    7432822,
    4852806,
    7211878,
    7668595,
    8127101,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    7733370,
    8391815,
    7274615,
    7996544,
    7864442,
    8389505,
    7471221,
    8324225,
    8783748,
    8915329,
    8456314,
    7080807,
    5710681,
    7825785,
    6912612,
    10865827,
    10801579,
    10407334,
    10210208,
    10407582,
    10934432,
    8829309,
    8171376,
    8698487,
    5146949,
    8303996,
    3825983,
    6975343,
    2949165,
    7411571,
    7405690,
    8652943,
    8323458,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    7799933,
    7608195,
    6559356,
    5770609,
    6886524,
    7276149,
    7932538,
    7801209,
    8064638,
    7998843,
    7802997,
    7148135,
    5511505,
    7761791,
    11521722,
    10804394,
    10018207,
    9952932,
    9755553,
    9689755,
    9821850,
    9427088,
    10348442,
    4361531,
    4887107,
    8505216,
    8371842,
    5473114,
    4740941,
    1966113,
    6033504,
    7603583,
    8257673,
    8454276,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8257917,
    8323197,
    7211641,
    4463210,
    3746156,
    4339062,
    4400749,
    6168434,
    6361963,
    6625134,
    6032998,
    5967972,
    5050711,
    5321567,
    7500165,
    11257794,
    10078901,
    9491379,
    9559221,
    9624242,
    1004843,
    12546,
    3768653,
    4690005,
    4427085,
    9822109,
    7586685,
    6601332,
    6929019,
    5278297,
    4086339,
    1313307,
    5775708,
    7933050,
    9045384,
    8519808,
    8454528,
    8519810,
    8519810,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8257917,
    8323197,
    6753909,
    8024491,
    11653874,
    11194861,
    3230058,
    4011104,
    4862050,
    7033478,
    7034248,
    6574464,
    6117757,
    4744303,
    4157545,
    4029802,
    2585176,
    2454620,
    152119,
    875324,
    10019520,
    9293485,
    11526,
    9030812,
    9361310,
    9230744,
    9100952,
    6932866,
    6404984,
    7518591,
    3499069,
    6782324,
    2100009,
    6426976,
    7602288,
    8454526,
    8519810,
    8519810,
    8519810,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8257917,
    8323197,
    8323197,
    8257917,
    8323197,
    8454269,
    6557809,
    6977433,
    10610149,
    9232080,
    9955287,
    3765099,
    3630949,
    10605272,
    10672348,
    10279128,
    10017748,
    9890264,
    7590841,
    6934706,
    7066292,
    22589,
    9694416,
    9694666,
    10217415,
    10143924,
    8203,
    10343597,
    9557406,
    9297298,
    8707469,
    6865785,
    6602618,
    7258235,
    2716472,
    4752734,
    6323573,
    2229033,
    6953834,
    8061819,
    8716422,
    8650884,
    8519810,
    8519810,
    8519810,
    8519810,
    8519810,
    8519810,
    8519810,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8257917,
    8323197,
    8323197,
    8323197,
    8323197,
    8454269,
    6361711,
    6849177,
    9167568,
    3776894,
    8119997,
    9234628,
    9628621,
    8708814,
    8643793,
    3577214,
    3709311,
    3316606,
    8581843,
    6150582,
    5886640,
    7724738,
    8512454,
    8710853,
    7654315,
    9422002,
    8205,
    10934199,
    9621918,
    9692054,
    9431187,
    7259000,
    7324542,
    7061622,
    3245376,
    1468465,
    5738609,
    1252130,
    5054034,
    7538805,
    8650884,
    8519810,
    8519810,
    8519810,
    8519810,
    8519810,
    8519810,
    8519810,
    8519810,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8257917,
    8257915,
    8323195,
    8323195,
    8323195,
    8127099,
    5969517,
    6391193,
    1997414,
    8579783,
    9171915,
    9235399,
    8840902,
    8383698,
    3449226,
    4431753,
    3970173,
    4365701,
    8580046,
    7599311,
    5691828,
    6937275,
    6738354,
    7134649,
    6672301,
    7194028,
    5018234,
    9481,
    10014625,
    9757338,
    9298834,
    7783035,
    8111232,
    7060341,
    4165967,
    1600819,
    5083498,
    5666409,
    1771814,
    6754409,
    8192892,
    8454528,
    8519810,
    8519810,
    8519810,
    8519810,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8257917,
    8127099,
    8257915,
    8454267,
    8257915,
    7800187,
    5511533,
    4747395,
    8512205,
    8251332,
    7856055,
    9366215,
    9235147,
    3711882,
    2725246,
    3971715,
    3378806,
    8642246,
    9040084,
    7927763,
    6480317,
    6014633,
    7131317,
    6805686,
    6477237,
    6739128,
    3641206,
    7942,
    10737069,
    9362328,
    7981952,
    8044665,
    8438911,
    7520378,
    4100173,
    3968596,
    1729588,
    5080162,
    659990,
    6035549,
    7800948,
    8127099,
    8454528,
    8585347,
    8585347,
    8323199,
    8323199,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8127101,
    8061819,
    8127099,
    8323193,
    8192122,
    7473532,
    4856169,
    4024441,
    8380618,
    8384200,
    9041099,
    9826252,
    8837822,
    4102020,
    3774341,
    3842183,
    8711633,
    8580046,
    8843988,
    8647636,
    7264187,
    4824455,
    4034169,
    6998963,
    6278323,
    6740673,
    3841413,
    8460,
    10933428,
    7519104,
    7455096,
    8175994,
    8241787,
    5152089,
    4232275,
    4033874,
    2125366,
    4493142,
    6588015,
    3080239,
    7212393,
    7800437,
    8126588,
    8585347,
    8585347,
    8323199,
    8257917,
    8323199,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8127101,
    8061819,
    8127099,
    8061045,
    8324221,
    6818169,
    7356817,
    3163483,
    10018768,
    6933418,
    8316606,
    8905664,
    9233352,
    9429713,
    9496279,
    7987142,
    8712659,
    8120779,
    7262390,
    10151122,
    4289898,
    12047826,
    11786453,
    1070668,
    7458751,
    3383181,
    3906697,
    5343354,
    9739,
    7452546,
    7389049,
    7585138,
    4230978,
    4365140,
    3443532,
    4362324,
    2059053,
    4627283,
    5078356,
    2557219,
    6754913,
    7669362,
    7995516,
    8585348,
    8585348,
    8192124,
    8061306,
    8257917,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8127101,
    7930749,
    8061821,
    8650876,
    8127612,
    6556537,
    5841009,
    6902132,
    7373443,
    9689537,
    7722672,
    9368013,
    8840906,
    9299156,
    4430220,
    3577984,
    8316105,
    6671536,
    10281938,
    5331295,
    7557734,
    6105409,
    16773119,
    12310495,
    1070418,
    4101005,
    3310458,
    5409408,
    7174,
    1727789,
    5020249,
    4035139,
    4497743,
    3512398,
    3050313,
    4887898,
    2321194,
    4034878,
    5539922,
    2165273,
    6493531,
    7407728,
    7995516,
    8585350,
    8585348,
    8192124,
    8061306,
    8257917,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8257917,
    8127101,
    8061821,
    8127101,
    8126582,
    7538294,
    5838960,
    5646696,
    8079211,
    9205889,
    11132618,
    7590319,
    8580296,
    8776655,
    3904646,
    3509118,
    3314040,
    8841419,
    7064497,
    11263189,
    7951979,
    9911650,
    8655932,
    16769791,
    16645631,
    1461331,
    4822677,
    3968906,
    4490623,
    11035,
    1004082,
    4362589,
    3838539,
    3576905,
    3182411,
    4167511,
    2584884,
    4361031,
    4560452,
    5407055,
    2492191,
    6689633,
    7538546,
    7995516,
    8585348,
    8585348,
    8192124,
    8061306,
    8257917,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8126847,
    8061567,
    8126847,
    8257917,
    8061049,
    6753389,
    7033984,
    13878235,
    9194857,
    16772604,
    6195578,
    8774596,
    8843986,
    8777943,
    4364429,
    4363914,
    8381636,
    9171150,
    9233102,
    6916235,
    8734567,
    16766207,
    9766450,
    8591161,
    16775167,
    11262691,
    3641742,
    4170394,
    4231562,
    807241,
    4294525,
    743486,
    3641180,
    3904087,
    3967570,
    5347938,
    1795883,
    4229706,
    5084752,
    6060124,
    3604533,
    7406703,
    8523138,
    7929976,
    8323201,
    8323201,
    8257917,
    8127101,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8061567,
    8061567,
    8126847,
    8257663,
    8061308,
    6097510,
    5921397,
    16121599,
    5973049,
    16772604,
    5868410,
    7461048,
    8187598,
    8515800,
    8708564,
    8906197,
    9107156,
    8382663,
    7851708,
    6390661,
    6105411,
    16769279,
    15890839,
    13596045,
    16774399,
    11591400,
    4167316,
    2986889,
    4233874,
    2783862,
    4952980,
    4492935,
    21305,
    4363632,
    4360804,
    2189372,
    3901773,
    4821330,
    5079119,
    1052688,
    6360929,
    8324223,
    8456064,
    8192894,
    8257663,
    8257663,
    8127101,
    8127101,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8126849,
    8061569,
    8061567,
    8061567,
    8061048,
    7018614,
    5922433,
    10664128,
    5057852,
    4009523,
    4427640,
    6215860,
    6084535,
    5952183,
    6805697,
    6542526,
    5755059,
    6214326,
    6868408,
    5410440,
    3617852,
    5911099,
    11962760,
    10980490,
    12570840,
    5670799,
    5216409,
    4298900,
    3906195,
    3904655,
    4492429,
    4820880,
    4493968,
    284496,
    350025,
    3968878,
    4956514,
    5214291,
    6254685,
    2754341,
    7608180,
    8390017,
    8324223,
    8455810,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323201,
    8257667,
    8126851,
    7930751,
    8061567,
    8520321,
    7082872,
    3748707,
    5672,
    11577782,
    10857646,
    9094584,
    7458999,
    6607799,
    6412475,
    6148535,
    6410938,
    6280122,
    6870975,
    7328444,
    8505529,
    10138797,
    11515823,
    10332567,
    10006432,
    6062723,
    5934998,
    938580,
    4033931,
    3642253,
    3904655,
    5085335,
    5084055,
    4689814,
    4953500,
    4757654,
    612677,
    4296794,
    5867358,
    1640473,
    6693476,
    7210092,
    8192894,
    8455810,
    8192894,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323201,
    8323205,
    8257669,
    7930751,
    8061821,
    8126588,
    7015030,
    4794219,
    7436187,
    4896,
    2767681,
    11645372,
    11321538,
    4757123,
    6869942,
    7789762,
    1802086,
    6473389,
    7787451,
    7652269,
    8569003,
    9156004,
    10536885,
    3763289,
    1001530,
    8480,
    7457,
    4558478,
    3902345,
    2389106,
    4494482,
    4231310,
    4229511,
    1134415,
    1396817,
    5214610,
    4754563,
    1396787,
    531223,
    5710433,
    6948719,
    7931001,
    8257917,
    8257917,
    8257917,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8585351,
    8454279,
    8126847,
    8061821,
    8323712,
    7735934,
    5180003,
    4598373,
    7306132,
    15728639,
    3680572,
    3617600,
    9419956,
    9225654,
    10009524,
    10664887,
    10138797,
    5729637,
    3819326,
    1056274,
    136969,
    6926,
    13762559,
    2650218,
    5279374,
    5344142,
    5083539,
    4690064,
    743767,
    4033931,
    4692372,
    4690830,
    1726034,
    1593934,
    1266514,
    5477520,
    5211513,
    3095882,
    5906795,
    6619502,
    7931003,
    8257917,
    8257917,
    8257917,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454275,
    8650889,
    8650887,
    8454271,
    8257915,
    7733372,
    8325509,
    7932538,
    6558313,
    4861018,
    7961746,
    7176332,
    5268584,
    3159610,
    4532278,
    7347772,
    9117506,
    7934253,
    8329520,
    8133163,
    7217451,
    5451059,
    3619907,
    3960697,
    4295059,
    4688529,
    5477016,
    5869207,
    936783,
    4100494,
    4102289,
    4034953,
    5414807,
    4755591,
    1070670,
    545356,
    4492168,
    5214092,
    6324366,
    5059172,
    6165863,
    7538805,
    8257917,
    8257917,
    8257917,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8650887,
    8650885,
    8585341,
    8323197,
    7471225,
    7864444,
    8650876,
    7799663,
    6955628,
    2360630,
    856883,
    7306898,
    7762305,
    7753312,
    7082547,
    11681635,
    14970770,
    14971533,
    14249345,
    13137794,
    8542816,
    7698560,
    5538961,
    4491929,
    5544356,
    8747,
    10548,
    4819086,
    3706761,
    4168849,
    4034181,
    4427910,
    2717806,
    4494216,
    4625034,
    4690316,
    5018516,
    5538961,
    3422296,
    4528470,
    7211891,
    8257917,
    8257917,
    8257917,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454273,
    8454273,
    8454269,
    8323197,
    8061056,
    8192128,
    8454270,
    8388730,
    8063352,
    6688366,
    5249644,
    1114167,
    3100,
    7046790,
    7240828,
    7895421,
    8417920,
    8614268,
    9075836,
    8881276,
    7570293,
    6720126,
    10024,
    9516,
    9009,
    4885142,
    4164754,
    3246214,
    2062192,
    3574659,
    4427140,
    611401,
    4167302,
    4101255,
    4558474,
    806992,
    4360331,
    4949137,
    6586521,
    1836862,
    6753907,
    8257917,
    8257917,
    8257917,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323199,
    8192126,
    8192128,
    8454270,
    8585342,
    7995507,
    8127614,
    6490230,
    5450870,
    6390420,
    10781,
    12317,
    7953,
    8738,
    9766,
    7958,
    8205,
    9485,
    7948,
    4754565,
    4886674,
    4426386,
    4165013,
    3510161,
    3445392,
    21582,
    4296072,
    5148298,
    12072,
    3576197,
    4233872,
    1136727,
    1397847,
    1003862,
    4488584,
    6458012,
    1511232,
    6688627,
    8257917,
    8257917,
    8257917,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8192126,
    8192126,
    8454270,
    8585342,
    8650878,
    7602293,
    7539838,
    9199275,
    9354442,
    6603440,
    7064758,
    4167302,
    938317,
    5409928,
    5608325,
    5083775,
    4758406,
    3640445,
    4887439,
    20044,
    7066574,
    6475466,
    3643798,
    3772558,
    4296333,
    1135443,
    5658,
    4949641,
    4168597,
    2919046,
    1004375,
    1067088,
    1199186,
    5473934,
    6062475,
    655658,
    6688625,
    8257917,
    8257917,
    8257917,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8192126,
    8192126,
    8454270,
    8454270,
    9046406,
    7929976,
    7997309,
    5512300,
    4222334,
    3446405,
    6737592,
    6932918,
    3967620,
    872270,
    12069,
    4686971,
    5081225,
    4556168,
    413004,
    4364177,
    3382931,
    6278595,
    7328460,
    3706765,
    4492429,
    1659223,
    6953,
    6130067,
    4627353,
    3971734,
    1071965,
    542285,
    1463127,
    5802386,
    6322567,
    2231609,
    6884975,
    8257917,
    8257917,
    8257917,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8454271,
    8585343,
    8519806,
    8257660,
    8324221,
    6035308,
    4614012,
    3642244,
    6473651,
    6999484,
    4231821,
    5083024,
    6460048,
    268580,
    1642038,
    855348,
    1463125,
    4365199,
    3640708,
    3773323,
    7393991,
    4300183,
    3702402,
    1656658,
    267563,
    6782866,
    4622988,
    4102291,
    4101007,
    613209,
    4756373,
    5342096,
    987951,
    4330575,
    7211889,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8454271,
    8585343,
    8650878,
    8519806,
    8454780,
    6558572,
    6977683,
    8833988,
    7391159,
    7590337,
    8049614,
    4426125,
    6390409,
    1445161,
    5380700,
    4662368,
    5737876,
    7260856,
    4362630,
    4231560,
    6670780,
    3640969,
    5736340,
    3425375,
    3221836,
    789543,
    3630183,
    5149321,
    2846827,
    4951437,
    3172980,
    6783132,
    2360632,
    5901916,
    7735157,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8454271,
    8585343,
    8716414,
    8650878,
    8454780,
    6885740,
    4140371,
    4877168,
    9226947,
    4495500,
    7130311,
    4690326,
    6518147,
    1900582,
    6100072,
    4988519,
    4947590,
    7524796,
    7324851,
    7852223,
    6408376,
    4756112,
    987438,
    5056342,
    5318235,
    4598864,
    12175300,
    2245171,
    12441300,
    2899017,
    12962282,
    4663905,
    6097760,
    7537258,
    8127097,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8454271,
    8585343,
    8716418,
    8716416,
    8454780,
    7277936,
    5646687,
    16709887,
    2835021,
    14942207,
    1265496,
    5931668,
    1837616,
    5511514,
    6886774,
    5052779,
    2575197,
    8177339,
    5148548,
    8832443,
    5149582,
    6588054,
    2228271,
    6362717,
    6164318,
    5509716,
    2294560,
    1771032,
    2295589,
    2424879,
    3080254,
    6100072,
    7932018,
    8782714,
    8454267,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8454271,
    8585345,
    8716424,
    8650888,
    8323712,
    7473782,
    6164833,
    3145782,
    1638434,
    2165036,
    1376806,
    2622775,
    6231912,
    6950772,
    6556791,
    6038392,
    16120575,
    2244682,
    15990783,
    3226437,
    16118783,
    2295607,
    6100322,
    7211630,
    7734390,
    7734390,
    7146348,
    6950248,
    7015532,
    7146096,
    7211380,
    7538294,
    8061306,
    8388732,
    8323197,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8454271,
    8585345,
    8716424,
    8650888,
    8323712,
    7800696,
    7343727,
    6623074,
    6164568,
    6231126,
    6361431,
    6687584,
    7867002,
    7603585,
    7080321,
    6099318,
    2687044,
    2032949,
    2097195,
    2949168,
    3539001,
    6362213,
    7146350,
    7865208,
    8388736,
    8585346,
    8388736,
    8257662,
    8257662,
    8257662,
    8257662,
    8257662,
    8257662,
    8257662,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8454271,
    8454271,
    8650880,
    8650880,
    8454780,
    8193144,
    7603055,
    7801200,
    7736942,
    7670382,
    8325496,
    8521857,
    8061058,
    8127112,
    7405698,
    7604100,
    7277436,
    7475579,
    7277686,
    7276919,
    7341429,
    7669112,
    7865210,
    8061308,
    8257662,
    8257662,
    8257662,
    8257660,
    8257662,
    8257662,
    8257662,
    8257662,
    8257662,
    8257662,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8257663,
    8323199,
    8323199,
    8454269,
    8650876,
    8520060,
    8520060,
    8454778,
    8718207,
    8258167,
    8061045,
    8323449,
    8126584,
    8716421,
    7995519,
    8389001,
    7995524,
    8323206,
    8061054,
    8061054,
    8192129,
    8783498,
    8061052,
    8389251,
    8192126,
    8192126,
    8192126,
    8192124,
    8257660,
    8257660,
    8257662,
    8257662,
    8257662,
    8257662,
    8257662,
    8257662,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8454269,
    8520060,
    8520060,
    8520060,
    8650878,
    8650878,
    8716416,
    8716416,
    8650880,
    8257665,
    8126849,
    8323199,
    8519806,
    8388732,
    8388734,
    8257664,
    8192126,
    8127097,
    8127351,
    8127097,
    8258169,
    8257915,
    8257917,
    8257663,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323197,
    8323197,
    8519808,
    8519808,
    8519808,
    8650880,
    8650882,
    8716418,
    8716418,
    8519810,
    8061569,
    8061567,
    8257917,
    8454269,
    8388732,
    8257660,
    8061054,
    8061308,
    8258167,
    8323701,
    8323701,
    8323447,
    8323195,
    8257917,
    8257917,
    8257663,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454271,
    8454273,
    8519814,
    8519816,
    8519814,
    8454276,
    8323458,
    8323458,
    8192640,
    8192640,
    8127101,
    8257917,
    8257665,
    8257667,
    8061058,
    7930240,
    7734140,
    7930490,
    8650873,
    8978553,
    8847481,
    8650875,
    8454267,
    8323197,
    8257917,
    8257917,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454271,
    8454273,
    8519814,
    8519816,
    8454278,
    8323460,
    8192642,
    8127360,
    8127360,
    8127614,
    8257917,
    8323197,
    8257665,
    8257667,
    8061058,
    7864704,
    7734140,
    8061308,
    8781949,
    8978557,
    8847485,
    8781949,
    8585341,
    8323197,
    8257917,
    8257917,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454274,
    8454274,
    8454274,
    8454274,
    8323712,
    8323712,
    8323712,
    8323712,
    8454528,
    8454528,
    8454528,
    8454274,
    8257665,
    8257663,
    8126847,
    8257663,
    8454271,
    8585343,
    8585343,
    8454271,
    8454271,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8454528,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199,
    8323199
  };

  always_ff @(posedge clk) begin
    if (!rst_n) begin
      o_rd_data <= '0;
    end else begin
      o_rd_data[0] <= bulbasaur_rom_buf[i_rd_addr];
      o_rd_data[1] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2];
    end
  end
endmodule
