module bulbasaur_rom_new #(
    parameter hpixel_p = 64,
    parameter vpixel_p = 64,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

    // Clock and reset
    input logic clk,
    input logic rst_n,

    /* Pixel read interface */
    input logic [addr_width_p-1:0] i_rd_addr,
    output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
    );


        logic [3*bpp_p-1:0] rd_data_0;
        logic [3*bpp_p-1:0] rd_data_1;

    always_ff @(posedge clk) begin
        case (i_rd_addr)
		12'd0000: rd_data_0 <= 24'h810081;
		12'd0001: rd_data_0 <= 24'h810081;
		12'd0002: rd_data_0 <= 24'h810081;
		12'd0003: rd_data_0 <= 24'h810081;
		12'd0004: rd_data_0 <= 24'h810081;
		12'd0005: rd_data_0 <= 24'h810081;
		12'd0006: rd_data_0 <= 24'h81007f;
		12'd0007: rd_data_0 <= 24'h81007f;
		12'd0008: rd_data_0 <= 24'h81007f;
		12'd0009: rd_data_0 <= 24'h81007f;
		12'd0010: rd_data_0 <= 24'h81007d;
		12'd0011: rd_data_0 <= 24'h81007d;
		12'd0012: rd_data_0 <= 24'h81007d;
		12'd0013: rd_data_0 <= 24'h81007d;
		12'd0014: rd_data_0 <= 24'h81007d;
		12'd0015: rd_data_0 <= 24'h81007d;
		12'd0016: rd_data_0 <= 24'h7f007f;
		12'd0017: rd_data_0 <= 24'h7f007f;
		12'd0018: rd_data_0 <= 24'h7f007f;
		12'd0019: rd_data_0 <= 24'h7f007f;
		12'd0020: rd_data_0 <= 24'h7f007f;
		12'd0021: rd_data_0 <= 24'h7f007f;
		12'd0022: rd_data_0 <= 24'h7f007f;
		12'd0023: rd_data_0 <= 24'h7f007f;
		12'd0024: rd_data_0 <= 24'h7f007f;
		12'd0025: rd_data_0 <= 24'h7f007f;
		12'd0026: rd_data_0 <= 24'h7f007f;
		12'd0027: rd_data_0 <= 24'h7f007f;
		12'd0028: rd_data_0 <= 24'h7f007f;
		12'd0029: rd_data_0 <= 24'h7f007f;
		12'd0030: rd_data_0 <= 24'h7f007f;
		12'd0031: rd_data_0 <= 24'h7f007f;
		12'd0032: rd_data_0 <= 24'h7f007f;
		12'd0033: rd_data_0 <= 24'h7f007f;
		12'd0034: rd_data_0 <= 24'h7f007f;
		12'd0035: rd_data_0 <= 24'h7f007f;
		12'd0036: rd_data_0 <= 24'h7f007f;
		12'd0037: rd_data_0 <= 24'h7f007f;
		12'd0038: rd_data_0 <= 24'h7f007f;
		12'd0039: rd_data_0 <= 24'h7f007f;
		12'd0040: rd_data_0 <= 24'h7f007f;
		12'd0041: rd_data_0 <= 24'h7f007f;
		12'd0042: rd_data_0 <= 24'h7f007f;
		12'd0043: rd_data_0 <= 24'h7f007f;
		12'd0044: rd_data_0 <= 24'h7f007f;
		12'd0045: rd_data_0 <= 24'h7f007f;
		12'd0046: rd_data_0 <= 24'h7f007f;
		12'd0047: rd_data_0 <= 24'h7f007f;
		12'd0048: rd_data_0 <= 24'h7f007f;
		12'd0049: rd_data_0 <= 24'h7f007f;
		12'd0050: rd_data_0 <= 24'h7f007f;
		12'd0051: rd_data_0 <= 24'h7f007f;
		12'd0052: rd_data_0 <= 24'h7f007f;
		12'd0053: rd_data_0 <= 24'h7f007f;
		12'd0054: rd_data_0 <= 24'h7f007f;
		12'd0055: rd_data_0 <= 24'h7f007f;
		12'd0056: rd_data_0 <= 24'h7f007f;
		12'd0057: rd_data_0 <= 24'h7f007f;
		12'd0058: rd_data_0 <= 24'h7f007f;
		12'd0059: rd_data_0 <= 24'h7f007f;
		12'd0060: rd_data_0 <= 24'h7f007f;
		12'd0061: rd_data_0 <= 24'h7f007f;
		12'd0062: rd_data_0 <= 24'h7f007f;
		12'd0063: rd_data_0 <= 24'h7f007f;
		12'd0064: rd_data_0 <= 24'h810081;
		12'd0065: rd_data_0 <= 24'h810081;
		12'd0066: rd_data_0 <= 24'h810081;
		12'd0067: rd_data_0 <= 24'h810081;
		12'd0068: rd_data_0 <= 24'h810081;
		12'd0069: rd_data_0 <= 24'h810081;
		12'd0070: rd_data_0 <= 24'h81007f;
		12'd0071: rd_data_0 <= 24'h81007f;
		12'd0072: rd_data_0 <= 24'h81007f;
		12'd0073: rd_data_0 <= 24'h81007f;
		12'd0074: rd_data_0 <= 24'h81007d;
		12'd0075: rd_data_0 <= 24'h81007d;
		12'd0076: rd_data_0 <= 24'h81007d;
		12'd0077: rd_data_0 <= 24'h81007d;
		12'd0078: rd_data_0 <= 24'h81007d;
		12'd0079: rd_data_0 <= 24'h81007d;
		12'd0080: rd_data_0 <= 24'h7f007f;
		12'd0081: rd_data_0 <= 24'h7f007f;
		12'd0082: rd_data_0 <= 24'h7f007f;
		12'd0083: rd_data_0 <= 24'h7f007f;
		12'd0084: rd_data_0 <= 24'h7f007f;
		12'd0085: rd_data_0 <= 24'h7f007f;
		12'd0086: rd_data_0 <= 24'h7f007f;
		12'd0087: rd_data_0 <= 24'h7f007f;
		12'd0088: rd_data_0 <= 24'h7f007f;
		12'd0089: rd_data_0 <= 24'h7f007f;
		12'd0090: rd_data_0 <= 24'h7f007f;
		12'd0091: rd_data_0 <= 24'h7f007f;
		12'd0092: rd_data_0 <= 24'h7f007f;
		12'd0093: rd_data_0 <= 24'h7f007f;
		12'd0094: rd_data_0 <= 24'h7f007f;
		12'd0095: rd_data_0 <= 24'h7f007f;
		12'd0096: rd_data_0 <= 24'h7f007f;
		12'd0097: rd_data_0 <= 24'h7f007f;
		12'd0098: rd_data_0 <= 24'h7f007f;
		12'd0099: rd_data_0 <= 24'h7f007f;
		12'd0100: rd_data_0 <= 24'h7f007f;
		12'd0101: rd_data_0 <= 24'h7f007f;
		12'd0102: rd_data_0 <= 24'h7f007f;
		12'd0103: rd_data_0 <= 24'h7f007f;
		12'd0104: rd_data_0 <= 24'h7f007f;
		12'd0105: rd_data_0 <= 24'h7f007f;
		12'd0106: rd_data_0 <= 24'h7f007f;
		12'd0107: rd_data_0 <= 24'h7f007f;
		12'd0108: rd_data_0 <= 24'h7f007f;
		12'd0109: rd_data_0 <= 24'h7f007f;
		12'd0110: rd_data_0 <= 24'h7f007f;
		12'd0111: rd_data_0 <= 24'h7f007f;
		12'd0112: rd_data_0 <= 24'h7f007f;
		12'd0113: rd_data_0 <= 24'h7f007f;
		12'd0114: rd_data_0 <= 24'h7f007f;
		12'd0115: rd_data_0 <= 24'h7f007f;
		12'd0116: rd_data_0 <= 24'h7f007f;
		12'd0117: rd_data_0 <= 24'h7f007f;
		12'd0118: rd_data_0 <= 24'h7f007f;
		12'd0119: rd_data_0 <= 24'h7f007f;
		12'd0120: rd_data_0 <= 24'h7f007f;
		12'd0121: rd_data_0 <= 24'h7f007f;
		12'd0122: rd_data_0 <= 24'h7f007f;
		12'd0123: rd_data_0 <= 24'h7f007f;
		12'd0124: rd_data_0 <= 24'h7f007f;
		12'd0125: rd_data_0 <= 24'h7f007f;
		12'd0126: rd_data_0 <= 24'h7f007f;
		12'd0127: rd_data_0 <= 24'h7f007f;
		12'd0128: rd_data_0 <= 24'h810081;
		12'd0129: rd_data_0 <= 24'h810081;
		12'd0130: rd_data_0 <= 24'h810081;
		12'd0131: rd_data_0 <= 24'h810081;
		12'd0132: rd_data_0 <= 24'h810081;
		12'd0133: rd_data_0 <= 24'h810081;
		12'd0134: rd_data_0 <= 24'h81007f;
		12'd0135: rd_data_0 <= 24'h81007f;
		12'd0136: rd_data_0 <= 24'h81007f;
		12'd0137: rd_data_0 <= 24'h81007f;
		12'd0138: rd_data_0 <= 24'h81007d;
		12'd0139: rd_data_0 <= 24'h81007d;
		12'd0140: rd_data_0 <= 24'h81007d;
		12'd0141: rd_data_0 <= 24'h81007d;
		12'd0142: rd_data_0 <= 24'h81007d;
		12'd0143: rd_data_0 <= 24'h81007d;
		12'd0144: rd_data_0 <= 24'h7f007f;
		12'd0145: rd_data_0 <= 24'h7f007f;
		12'd0146: rd_data_0 <= 24'h7f007f;
		12'd0147: rd_data_0 <= 24'h7f007f;
		12'd0148: rd_data_0 <= 24'h7f007f;
		12'd0149: rd_data_0 <= 24'h7f007f;
		12'd0150: rd_data_0 <= 24'h7f007f;
		12'd0151: rd_data_0 <= 24'h7f007f;
		12'd0152: rd_data_0 <= 24'h7f007f;
		12'd0153: rd_data_0 <= 24'h7f007f;
		12'd0154: rd_data_0 <= 24'h7f007f;
		12'd0155: rd_data_0 <= 24'h7f007f;
		12'd0156: rd_data_0 <= 24'h7f007f;
		12'd0157: rd_data_0 <= 24'h7f007f;
		12'd0158: rd_data_0 <= 24'h7f007f;
		12'd0159: rd_data_0 <= 24'h7f007f;
		12'd0160: rd_data_0 <= 24'h7f007f;
		12'd0161: rd_data_0 <= 24'h7f007f;
		12'd0162: rd_data_0 <= 24'h7f007f;
		12'd0163: rd_data_0 <= 24'h7f007f;
		12'd0164: rd_data_0 <= 24'h7f007f;
		12'd0165: rd_data_0 <= 24'h7f007f;
		12'd0166: rd_data_0 <= 24'h7f007f;
		12'd0167: rd_data_0 <= 24'h7f007f;
		12'd0168: rd_data_0 <= 24'h7f007f;
		12'd0169: rd_data_0 <= 24'h7f007f;
		12'd0170: rd_data_0 <= 24'h7f007f;
		12'd0171: rd_data_0 <= 24'h7f007f;
		12'd0172: rd_data_0 <= 24'h7f007f;
		12'd0173: rd_data_0 <= 24'h7f007f;
		12'd0174: rd_data_0 <= 24'h7f007f;
		12'd0175: rd_data_0 <= 24'h7f007f;
		12'd0176: rd_data_0 <= 24'h7f007f;
		12'd0177: rd_data_0 <= 24'h7f007f;
		12'd0178: rd_data_0 <= 24'h7f007f;
		12'd0179: rd_data_0 <= 24'h7f007f;
		12'd0180: rd_data_0 <= 24'h7f007f;
		12'd0181: rd_data_0 <= 24'h7f007f;
		12'd0182: rd_data_0 <= 24'h7f007f;
		12'd0183: rd_data_0 <= 24'h7f007f;
		12'd0184: rd_data_0 <= 24'h7f007f;
		12'd0185: rd_data_0 <= 24'h7f007f;
		12'd0186: rd_data_0 <= 24'h7f007f;
		12'd0187: rd_data_0 <= 24'h7f007f;
		12'd0188: rd_data_0 <= 24'h7f007f;
		12'd0189: rd_data_0 <= 24'h7f007f;
		12'd0190: rd_data_0 <= 24'h7f007f;
		12'd0191: rd_data_0 <= 24'h7f007f;
		12'd0192: rd_data_0 <= 24'h810081;
		12'd0193: rd_data_0 <= 24'h810081;
		12'd0194: rd_data_0 <= 24'h810081;
		12'd0195: rd_data_0 <= 24'h810081;
		12'd0196: rd_data_0 <= 24'h810081;
		12'd0197: rd_data_0 <= 24'h810081;
		12'd0198: rd_data_0 <= 24'h81007f;
		12'd0199: rd_data_0 <= 24'h81007f;
		12'd0200: rd_data_0 <= 24'h81007f;
		12'd0201: rd_data_0 <= 24'h81007f;
		12'd0202: rd_data_0 <= 24'h81007d;
		12'd0203: rd_data_0 <= 24'h81007d;
		12'd0204: rd_data_0 <= 24'h81007d;
		12'd0205: rd_data_0 <= 24'h81007d;
		12'd0206: rd_data_0 <= 24'h81007d;
		12'd0207: rd_data_0 <= 24'h81007d;
		12'd0208: rd_data_0 <= 24'h7f007f;
		12'd0209: rd_data_0 <= 24'h7f007f;
		12'd0210: rd_data_0 <= 24'h7f007f;
		12'd0211: rd_data_0 <= 24'h7f007f;
		12'd0212: rd_data_0 <= 24'h7f007f;
		12'd0213: rd_data_0 <= 24'h7f007f;
		12'd0214: rd_data_0 <= 24'h7f007f;
		12'd0215: rd_data_0 <= 24'h7f007f;
		12'd0216: rd_data_0 <= 24'h7f007f;
		12'd0217: rd_data_0 <= 24'h7f007f;
		12'd0218: rd_data_0 <= 24'h7f007f;
		12'd0219: rd_data_0 <= 24'h7f007f;
		12'd0220: rd_data_0 <= 24'h7f007f;
		12'd0221: rd_data_0 <= 24'h7f007f;
		12'd0222: rd_data_0 <= 24'h7f007f;
		12'd0223: rd_data_0 <= 24'h7f007f;
		12'd0224: rd_data_0 <= 24'h7f007f;
		12'd0225: rd_data_0 <= 24'h7f007f;
		12'd0226: rd_data_0 <= 24'h7f007f;
		12'd0227: rd_data_0 <= 24'h7f007f;
		12'd0228: rd_data_0 <= 24'h7f007f;
		12'd0229: rd_data_0 <= 24'h7f007f;
		12'd0230: rd_data_0 <= 24'h7f007f;
		12'd0231: rd_data_0 <= 24'h7f007f;
		12'd0232: rd_data_0 <= 24'h7f007f;
		12'd0233: rd_data_0 <= 24'h7f007f;
		12'd0234: rd_data_0 <= 24'h7f007f;
		12'd0235: rd_data_0 <= 24'h7f007f;
		12'd0236: rd_data_0 <= 24'h7f007f;
		12'd0237: rd_data_0 <= 24'h7f007f;
		12'd0238: rd_data_0 <= 24'h7f007f;
		12'd0239: rd_data_0 <= 24'h7f007f;
		12'd0240: rd_data_0 <= 24'h7f007f;
		12'd0241: rd_data_0 <= 24'h7f007f;
		12'd0242: rd_data_0 <= 24'h7f007f;
		12'd0243: rd_data_0 <= 24'h7f007f;
		12'd0244: rd_data_0 <= 24'h7f007f;
		12'd0245: rd_data_0 <= 24'h7f007f;
		12'd0246: rd_data_0 <= 24'h7f007f;
		12'd0247: rd_data_0 <= 24'h7f007f;
		12'd0248: rd_data_0 <= 24'h7f007f;
		12'd0249: rd_data_0 <= 24'h7f007f;
		12'd0250: rd_data_0 <= 24'h7f007f;
		12'd0251: rd_data_0 <= 24'h7f007f;
		12'd0252: rd_data_0 <= 24'h7f007f;
		12'd0253: rd_data_0 <= 24'h7f007f;
		12'd0254: rd_data_0 <= 24'h7f007f;
		12'd0255: rd_data_0 <= 24'h7f007f;
		12'd0256: rd_data_0 <= 24'h810081;
		12'd0257: rd_data_0 <= 24'h810081;
		12'd0258: rd_data_0 <= 24'h810081;
		12'd0259: rd_data_0 <= 24'h810081;
		12'd0260: rd_data_0 <= 24'h810081;
		12'd0261: rd_data_0 <= 24'h810081;
		12'd0262: rd_data_0 <= 24'h81007f;
		12'd0263: rd_data_0 <= 24'h81007f;
		12'd0264: rd_data_0 <= 24'h81007f;
		12'd0265: rd_data_0 <= 24'h81007f;
		12'd0266: rd_data_0 <= 24'h81007d;
		12'd0267: rd_data_0 <= 24'h81007d;
		12'd0268: rd_data_0 <= 24'h81007f;
		12'd0269: rd_data_0 <= 24'h81007f;
		12'd0270: rd_data_0 <= 24'h81007f;
		12'd0271: rd_data_0 <= 24'h81007f;
		12'd0272: rd_data_0 <= 24'h7f007f;
		12'd0273: rd_data_0 <= 24'h7f007f;
		12'd0274: rd_data_0 <= 24'h7f007f;
		12'd0275: rd_data_0 <= 24'h7f007f;
		12'd0276: rd_data_0 <= 24'h7f007f;
		12'd0277: rd_data_0 <= 24'h7f007f;
		12'd0278: rd_data_0 <= 24'h7f007f;
		12'd0279: rd_data_0 <= 24'h7f007f;
		12'd0280: rd_data_0 <= 24'h7f007f;
		12'd0281: rd_data_0 <= 24'h7f007f;
		12'd0282: rd_data_0 <= 24'h7f007f;
		12'd0283: rd_data_0 <= 24'h7f007f;
		12'd0284: rd_data_0 <= 24'h7f007f;
		12'd0285: rd_data_0 <= 24'h7f007f;
		12'd0286: rd_data_0 <= 24'h7f007f;
		12'd0287: rd_data_0 <= 24'h7f007f;
		12'd0288: rd_data_0 <= 24'h7f007f;
		12'd0289: rd_data_0 <= 24'h7f007f;
		12'd0290: rd_data_0 <= 24'h7f007f;
		12'd0291: rd_data_0 <= 24'h7f007f;
		12'd0292: rd_data_0 <= 24'h7f007f;
		12'd0293: rd_data_0 <= 24'h7f007f;
		12'd0294: rd_data_0 <= 24'h7f007f;
		12'd0295: rd_data_0 <= 24'h7f007f;
		12'd0296: rd_data_0 <= 24'h7f007f;
		12'd0297: rd_data_0 <= 24'h7f007f;
		12'd0298: rd_data_0 <= 24'h7f007f;
		12'd0299: rd_data_0 <= 24'h7f007f;
		12'd0300: rd_data_0 <= 24'h7f007f;
		12'd0301: rd_data_0 <= 24'h7f007f;
		12'd0302: rd_data_0 <= 24'h7f007f;
		12'd0303: rd_data_0 <= 24'h7f007f;
		12'd0304: rd_data_0 <= 24'h7f007f;
		12'd0305: rd_data_0 <= 24'h7f007f;
		12'd0306: rd_data_0 <= 24'h7f007f;
		12'd0307: rd_data_0 <= 24'h7f007f;
		12'd0308: rd_data_0 <= 24'h7f007f;
		12'd0309: rd_data_0 <= 24'h7f007f;
		12'd0310: rd_data_0 <= 24'h7f007f;
		12'd0311: rd_data_0 <= 24'h7f007f;
		12'd0312: rd_data_0 <= 24'h7f007f;
		12'd0313: rd_data_0 <= 24'h7f007f;
		12'd0314: rd_data_0 <= 24'h7f007f;
		12'd0315: rd_data_0 <= 24'h7f007f;
		12'd0316: rd_data_0 <= 24'h7f007f;
		12'd0317: rd_data_0 <= 24'h7f007f;
		12'd0318: rd_data_0 <= 24'h7f007f;
		12'd0319: rd_data_0 <= 24'h7f007f;
		12'd0320: rd_data_0 <= 24'h810081;
		12'd0321: rd_data_0 <= 24'h810081;
		12'd0322: rd_data_0 <= 24'h810081;
		12'd0323: rd_data_0 <= 24'h810081;
		12'd0324: rd_data_0 <= 24'h810081;
		12'd0325: rd_data_0 <= 24'h810081;
		12'd0326: rd_data_0 <= 24'h81007f;
		12'd0327: rd_data_0 <= 24'h81007f;
		12'd0328: rd_data_0 <= 24'h81007f;
		12'd0329: rd_data_0 <= 24'h81007f;
		12'd0330: rd_data_0 <= 24'h81007d;
		12'd0331: rd_data_0 <= 24'h81007d;
		12'd0332: rd_data_0 <= 24'h81007f;
		12'd0333: rd_data_0 <= 24'h81007f;
		12'd0334: rd_data_0 <= 24'h81007f;
		12'd0335: rd_data_0 <= 24'h81007f;
		12'd0336: rd_data_0 <= 24'h7f007f;
		12'd0337: rd_data_0 <= 24'h7f007f;
		12'd0338: rd_data_0 <= 24'h7f007f;
		12'd0339: rd_data_0 <= 24'h7f007f;
		12'd0340: rd_data_0 <= 24'h7f007f;
		12'd0341: rd_data_0 <= 24'h7f007f;
		12'd0342: rd_data_0 <= 24'h7f007f;
		12'd0343: rd_data_0 <= 24'h7f007f;
		12'd0344: rd_data_0 <= 24'h7f007f;
		12'd0345: rd_data_0 <= 24'h7f007f;
		12'd0346: rd_data_0 <= 24'h7f007f;
		12'd0347: rd_data_0 <= 24'h7f007f;
		12'd0348: rd_data_0 <= 24'h7f007f;
		12'd0349: rd_data_0 <= 24'h7f007f;
		12'd0350: rd_data_0 <= 24'h7f007f;
		12'd0351: rd_data_0 <= 24'h7f007f;
		12'd0352: rd_data_0 <= 24'h7f007f;
		12'd0353: rd_data_0 <= 24'h7f007f;
		12'd0354: rd_data_0 <= 24'h7f007f;
		12'd0355: rd_data_0 <= 24'h7f007f;
		12'd0356: rd_data_0 <= 24'h7f007f;
		12'd0357: rd_data_0 <= 24'h7f007f;
		12'd0358: rd_data_0 <= 24'h7f007f;
		12'd0359: rd_data_0 <= 24'h7f007f;
		12'd0360: rd_data_0 <= 24'h7f007f;
		12'd0361: rd_data_0 <= 24'h7f007f;
		12'd0362: rd_data_0 <= 24'h7f007f;
		12'd0363: rd_data_0 <= 24'h7f007f;
		12'd0364: rd_data_0 <= 24'h7f007f;
		12'd0365: rd_data_0 <= 24'h7f007f;
		12'd0366: rd_data_0 <= 24'h7f007f;
		12'd0367: rd_data_0 <= 24'h7f007f;
		12'd0368: rd_data_0 <= 24'h7f007f;
		12'd0369: rd_data_0 <= 24'h7f007f;
		12'd0370: rd_data_0 <= 24'h7f007f;
		12'd0371: rd_data_0 <= 24'h7f007f;
		12'd0372: rd_data_0 <= 24'h7f007f;
		12'd0373: rd_data_0 <= 24'h7f007f;
		12'd0374: rd_data_0 <= 24'h7f007f;
		12'd0375: rd_data_0 <= 24'h7f007f;
		12'd0376: rd_data_0 <= 24'h7f007f;
		12'd0377: rd_data_0 <= 24'h7f007f;
		12'd0378: rd_data_0 <= 24'h7f007f;
		12'd0379: rd_data_0 <= 24'h7f007f;
		12'd0380: rd_data_0 <= 24'h7f007f;
		12'd0381: rd_data_0 <= 24'h7f007f;
		12'd0382: rd_data_0 <= 24'h7f007f;
		12'd0383: rd_data_0 <= 24'h7f007f;
		12'd0384: rd_data_0 <= 24'h81007f;
		12'd0385: rd_data_0 <= 24'h81007f;
		12'd0386: rd_data_0 <= 24'h81007f;
		12'd0387: rd_data_0 <= 24'h81007f;
		12'd0388: rd_data_0 <= 24'h810081;
		12'd0389: rd_data_0 <= 24'h810081;
		12'd0390: rd_data_0 <= 24'h81007f;
		12'd0391: rd_data_0 <= 24'h81007f;
		12'd0392: rd_data_0 <= 24'h7f007f;
		12'd0393: rd_data_0 <= 24'h7f007f;
		12'd0394: rd_data_0 <= 24'h7f007d;
		12'd0395: rd_data_0 <= 24'h7f007d;
		12'd0396: rd_data_0 <= 24'h7f007f;
		12'd0397: rd_data_0 <= 24'h7f007f;
		12'd0398: rd_data_0 <= 24'h7f007f;
		12'd0399: rd_data_0 <= 24'h7f007f;
		12'd0400: rd_data_0 <= 24'h7f007f;
		12'd0401: rd_data_0 <= 24'h7f007f;
		12'd0402: rd_data_0 <= 24'h7f007f;
		12'd0403: rd_data_0 <= 24'h7f007f;
		12'd0404: rd_data_0 <= 24'h7f007f;
		12'd0405: rd_data_0 <= 24'h7f007f;
		12'd0406: rd_data_0 <= 24'h7f007f;
		12'd0407: rd_data_0 <= 24'h7f007f;
		12'd0408: rd_data_0 <= 24'h7f007f;
		12'd0409: rd_data_0 <= 24'h7f007f;
		12'd0410: rd_data_0 <= 24'h7f007f;
		12'd0411: rd_data_0 <= 24'h7f007f;
		12'd0412: rd_data_0 <= 24'h7f007f;
		12'd0413: rd_data_0 <= 24'h7f007f;
		12'd0414: rd_data_0 <= 24'h7f007f;
		12'd0415: rd_data_0 <= 24'h7f007f;
		12'd0416: rd_data_0 <= 24'h7f007f;
		12'd0417: rd_data_0 <= 24'h7f007f;
		12'd0418: rd_data_0 <= 24'h7f007f;
		12'd0419: rd_data_0 <= 24'h7f007f;
		12'd0420: rd_data_0 <= 24'h7f007f;
		12'd0421: rd_data_0 <= 24'h7f007f;
		12'd0422: rd_data_0 <= 24'h7f007f;
		12'd0423: rd_data_0 <= 24'h7f007f;
		12'd0424: rd_data_0 <= 24'h7f007f;
		12'd0425: rd_data_0 <= 24'h7f007f;
		12'd0426: rd_data_0 <= 24'h7f007f;
		12'd0427: rd_data_0 <= 24'h7f007f;
		12'd0428: rd_data_0 <= 24'h7f007f;
		12'd0429: rd_data_0 <= 24'h7f007f;
		12'd0430: rd_data_0 <= 24'h7f007f;
		12'd0431: rd_data_0 <= 24'h7f007f;
		12'd0432: rd_data_0 <= 24'h7f007f;
		12'd0433: rd_data_0 <= 24'h7f007f;
		12'd0434: rd_data_0 <= 24'h7f007f;
		12'd0435: rd_data_0 <= 24'h7f007f;
		12'd0436: rd_data_0 <= 24'h7f007f;
		12'd0437: rd_data_0 <= 24'h7f007f;
		12'd0438: rd_data_0 <= 24'h7f007f;
		12'd0439: rd_data_0 <= 24'h7f007f;
		12'd0440: rd_data_0 <= 24'h7f007f;
		12'd0441: rd_data_0 <= 24'h7f007f;
		12'd0442: rd_data_0 <= 24'h7f007f;
		12'd0443: rd_data_0 <= 24'h7f007f;
		12'd0444: rd_data_0 <= 24'h7f007f;
		12'd0445: rd_data_0 <= 24'h7f007f;
		12'd0446: rd_data_0 <= 24'h7f007f;
		12'd0447: rd_data_0 <= 24'h7f007f;
		12'd0448: rd_data_0 <= 24'h81007f;
		12'd0449: rd_data_0 <= 24'h81007f;
		12'd0450: rd_data_0 <= 24'h81007f;
		12'd0451: rd_data_0 <= 24'h81007f;
		12'd0452: rd_data_0 <= 24'h810081;
		12'd0453: rd_data_0 <= 24'h810081;
		12'd0454: rd_data_0 <= 24'h81007f;
		12'd0455: rd_data_0 <= 24'h81007f;
		12'd0456: rd_data_0 <= 24'h7f007f;
		12'd0457: rd_data_0 <= 24'h7f007f;
		12'd0458: rd_data_0 <= 24'h7f007d;
		12'd0459: rd_data_0 <= 24'h7f007d;
		12'd0460: rd_data_0 <= 24'h7f007f;
		12'd0461: rd_data_0 <= 24'h7f007f;
		12'd0462: rd_data_0 <= 24'h7f007f;
		12'd0463: rd_data_0 <= 24'h7f007f;
		12'd0464: rd_data_0 <= 24'h7f007f;
		12'd0465: rd_data_0 <= 24'h7f007f;
		12'd0466: rd_data_0 <= 24'h7f007f;
		12'd0467: rd_data_0 <= 24'h7f007f;
		12'd0468: rd_data_0 <= 24'h7f007f;
		12'd0469: rd_data_0 <= 24'h7f007f;
		12'd0470: rd_data_0 <= 24'h7f007f;
		12'd0471: rd_data_0 <= 24'h7f007f;
		12'd0472: rd_data_0 <= 24'h7f007f;
		12'd0473: rd_data_0 <= 24'h7f007f;
		12'd0474: rd_data_0 <= 24'h7f007f;
		12'd0475: rd_data_0 <= 24'h7f007f;
		12'd0476: rd_data_0 <= 24'h7f007f;
		12'd0477: rd_data_0 <= 24'h7f007f;
		12'd0478: rd_data_0 <= 24'h7f007f;
		12'd0479: rd_data_0 <= 24'h7f007f;
		12'd0480: rd_data_0 <= 24'h7f007f;
		12'd0481: rd_data_0 <= 24'h7f007f;
		12'd0482: rd_data_0 <= 24'h7f007f;
		12'd0483: rd_data_0 <= 24'h7f007f;
		12'd0484: rd_data_0 <= 24'h7f007f;
		12'd0485: rd_data_0 <= 24'h7f007f;
		12'd0486: rd_data_0 <= 24'h7f007f;
		12'd0487: rd_data_0 <= 24'h7f007f;
		12'd0488: rd_data_0 <= 24'h7f007f;
		12'd0489: rd_data_0 <= 24'h7f007f;
		12'd0490: rd_data_0 <= 24'h7f007f;
		12'd0491: rd_data_0 <= 24'h7f007f;
		12'd0492: rd_data_0 <= 24'h7f007f;
		12'd0493: rd_data_0 <= 24'h7f007f;
		12'd0494: rd_data_0 <= 24'h7f007f;
		12'd0495: rd_data_0 <= 24'h7f007f;
		12'd0496: rd_data_0 <= 24'h7f007f;
		12'd0497: rd_data_0 <= 24'h7f007f;
		12'd0498: rd_data_0 <= 24'h7f007f;
		12'd0499: rd_data_0 <= 24'h7f007f;
		12'd0500: rd_data_0 <= 24'h7f007f;
		12'd0501: rd_data_0 <= 24'h7f007f;
		12'd0502: rd_data_0 <= 24'h7f007f;
		12'd0503: rd_data_0 <= 24'h7f007f;
		12'd0504: rd_data_0 <= 24'h7f007f;
		12'd0505: rd_data_0 <= 24'h7f007f;
		12'd0506: rd_data_0 <= 24'h7f007f;
		12'd0507: rd_data_0 <= 24'h7f007f;
		12'd0508: rd_data_0 <= 24'h7f007f;
		12'd0509: rd_data_0 <= 24'h7f007f;
		12'd0510: rd_data_0 <= 24'h7f007f;
		12'd0511: rd_data_0 <= 24'h7f007f;
		12'd0512: rd_data_0 <= 24'h81007f;
		12'd0513: rd_data_0 <= 24'h81007f;
		12'd0514: rd_data_0 <= 24'h81007f;
		12'd0515: rd_data_0 <= 24'h81007f;
		12'd0516: rd_data_0 <= 24'h81007f;
		12'd0517: rd_data_0 <= 24'h81007f;
		12'd0518: rd_data_0 <= 24'h7f007f;
		12'd0519: rd_data_0 <= 24'h7f007f;
		12'd0520: rd_data_0 <= 24'h7f007f;
		12'd0521: rd_data_0 <= 24'h7f007f;
		12'd0522: rd_data_0 <= 24'h7e007f;
		12'd0523: rd_data_0 <= 24'h7e007f;
		12'd0524: rd_data_0 <= 24'h7e007f;
		12'd0525: rd_data_0 <= 24'h7e007f;
		12'd0526: rd_data_0 <= 24'h7e007f;
		12'd0527: rd_data_0 <= 24'h7e007f;
		12'd0528: rd_data_0 <= 24'h7f007f;
		12'd0529: rd_data_0 <= 24'h7f007f;
		12'd0530: rd_data_0 <= 24'h7f007f;
		12'd0531: rd_data_0 <= 24'h7f007f;
		12'd0532: rd_data_0 <= 24'h7f007f;
		12'd0533: rd_data_0 <= 24'h7f007f;
		12'd0534: rd_data_0 <= 24'h7f007f;
		12'd0535: rd_data_0 <= 24'h7f007f;
		12'd0536: rd_data_0 <= 24'h7f007f;
		12'd0537: rd_data_0 <= 24'h7f007f;
		12'd0538: rd_data_0 <= 24'h7f007f;
		12'd0539: rd_data_0 <= 24'h7f007f;
		12'd0540: rd_data_0 <= 24'h7f007f;
		12'd0541: rd_data_0 <= 24'h7f007f;
		12'd0542: rd_data_0 <= 24'h7f007f;
		12'd0543: rd_data_0 <= 24'h7f007f;
		12'd0544: rd_data_0 <= 24'h7f007f;
		12'd0545: rd_data_0 <= 24'h7f007f;
		12'd0546: rd_data_0 <= 24'h7f007f;
		12'd0547: rd_data_0 <= 24'h7f007f;
		12'd0548: rd_data_0 <= 24'h7f007f;
		12'd0549: rd_data_0 <= 24'h7f007f;
		12'd0550: rd_data_0 <= 24'h7f007f;
		12'd0551: rd_data_0 <= 24'h7f007f;
		12'd0552: rd_data_0 <= 24'h7f007f;
		12'd0553: rd_data_0 <= 24'h7f007f;
		12'd0554: rd_data_0 <= 24'h7f007f;
		12'd0555: rd_data_0 <= 24'h7f007f;
		12'd0556: rd_data_0 <= 24'h7f007f;
		12'd0557: rd_data_0 <= 24'h7f007f;
		12'd0558: rd_data_0 <= 24'h7f007f;
		12'd0559: rd_data_0 <= 24'h7f007f;
		12'd0560: rd_data_0 <= 24'h7f007f;
		12'd0561: rd_data_0 <= 24'h7f007f;
		12'd0562: rd_data_0 <= 24'h7f007f;
		12'd0563: rd_data_0 <= 24'h7f007f;
		12'd0564: rd_data_0 <= 24'h7f007f;
		12'd0565: rd_data_0 <= 24'h7f007f;
		12'd0566: rd_data_0 <= 24'h7f007f;
		12'd0567: rd_data_0 <= 24'h7f007f;
		12'd0568: rd_data_0 <= 24'h7f007f;
		12'd0569: rd_data_0 <= 24'h7f007f;
		12'd0570: rd_data_0 <= 24'h7f007f;
		12'd0571: rd_data_0 <= 24'h7f007f;
		12'd0572: rd_data_0 <= 24'h7f007f;
		12'd0573: rd_data_0 <= 24'h7f007f;
		12'd0574: rd_data_0 <= 24'h7f007f;
		12'd0575: rd_data_0 <= 24'h7f007f;
		12'd0576: rd_data_0 <= 24'h81007f;
		12'd0577: rd_data_0 <= 24'h81007f;
		12'd0578: rd_data_0 <= 24'h81007f;
		12'd0579: rd_data_0 <= 24'h81007f;
		12'd0580: rd_data_0 <= 24'h81007f;
		12'd0581: rd_data_0 <= 24'h81007f;
		12'd0582: rd_data_0 <= 24'h7f007f;
		12'd0583: rd_data_0 <= 24'h7f007f;
		12'd0584: rd_data_0 <= 24'h7f007f;
		12'd0585: rd_data_0 <= 24'h7f007f;
		12'd0586: rd_data_0 <= 24'h7e007f;
		12'd0587: rd_data_0 <= 24'h7e007f;
		12'd0588: rd_data_0 <= 24'h7e007f;
		12'd0589: rd_data_0 <= 24'h7e007f;
		12'd0590: rd_data_0 <= 24'h7e007f;
		12'd0591: rd_data_0 <= 24'h7e007f;
		12'd0592: rd_data_0 <= 24'h7f007f;
		12'd0593: rd_data_0 <= 24'h7f007f;
		12'd0594: rd_data_0 <= 24'h7f007f;
		12'd0595: rd_data_0 <= 24'h7f007f;
		12'd0596: rd_data_0 <= 24'h7f007f;
		12'd0597: rd_data_0 <= 24'h7f007f;
		12'd0598: rd_data_0 <= 24'h7f007f;
		12'd0599: rd_data_0 <= 24'h7f007f;
		12'd0600: rd_data_0 <= 24'h7f007f;
		12'd0601: rd_data_0 <= 24'h7f007f;
		12'd0602: rd_data_0 <= 24'h7f007f;
		12'd0603: rd_data_0 <= 24'h7f007f;
		12'd0604: rd_data_0 <= 24'h7f007f;
		12'd0605: rd_data_0 <= 24'h7f007f;
		12'd0606: rd_data_0 <= 24'h7f007f;
		12'd0607: rd_data_0 <= 24'h7f007f;
		12'd0608: rd_data_0 <= 24'h7f007f;
		12'd0609: rd_data_0 <= 24'h7f007f;
		12'd0610: rd_data_0 <= 24'h7f007f;
		12'd0611: rd_data_0 <= 24'h7f007f;
		12'd0612: rd_data_0 <= 24'h7f007f;
		12'd0613: rd_data_0 <= 24'h7f007f;
		12'd0614: rd_data_0 <= 24'h7f007f;
		12'd0615: rd_data_0 <= 24'h7f007f;
		12'd0616: rd_data_0 <= 24'h7f007f;
		12'd0617: rd_data_0 <= 24'h7f007f;
		12'd0618: rd_data_0 <= 24'h7f007f;
		12'd0619: rd_data_0 <= 24'h7f007f;
		12'd0620: rd_data_0 <= 24'h7f007f;
		12'd0621: rd_data_0 <= 24'h7f007f;
		12'd0622: rd_data_0 <= 24'h7f007f;
		12'd0623: rd_data_0 <= 24'h7f007f;
		12'd0624: rd_data_0 <= 24'h7f007f;
		12'd0625: rd_data_0 <= 24'h7f007f;
		12'd0626: rd_data_0 <= 24'h7f007f;
		12'd0627: rd_data_0 <= 24'h7f007f;
		12'd0628: rd_data_0 <= 24'h7f007f;
		12'd0629: rd_data_0 <= 24'h7f007f;
		12'd0630: rd_data_0 <= 24'h7f007f;
		12'd0631: rd_data_0 <= 24'h7f007f;
		12'd0632: rd_data_0 <= 24'h7f007f;
		12'd0633: rd_data_0 <= 24'h7f007f;
		12'd0634: rd_data_0 <= 24'h7f007f;
		12'd0635: rd_data_0 <= 24'h7f007f;
		12'd0636: rd_data_0 <= 24'h7f007f;
		12'd0637: rd_data_0 <= 24'h7f007f;
		12'd0638: rd_data_0 <= 24'h7f007f;
		12'd0639: rd_data_0 <= 24'h7f007f;
		12'd0640: rd_data_0 <= 24'h81007d;
		12'd0641: rd_data_0 <= 24'h81007d;
		12'd0642: rd_data_0 <= 24'h81007d;
		12'd0643: rd_data_0 <= 24'h81007d;
		12'd0644: rd_data_0 <= 24'h81007f;
		12'd0645: rd_data_0 <= 24'h81007f;
		12'd0646: rd_data_0 <= 24'h7f007f;
		12'd0647: rd_data_0 <= 24'h7f007f;
		12'd0648: rd_data_0 <= 24'h7e007f;
		12'd0649: rd_data_0 <= 24'h7e007f;
		12'd0650: rd_data_0 <= 24'h7e007f;
		12'd0651: rd_data_0 <= 24'h7c017f;
		12'd0652: rd_data_0 <= 24'h7e007f;
		12'd0653: rd_data_0 <= 24'h7e007f;
		12'd0654: rd_data_0 <= 24'h7e007f;
		12'd0655: rd_data_0 <= 24'h7e007f;
		12'd0656: rd_data_0 <= 24'h7e007f;
		12'd0657: rd_data_0 <= 24'h7e007f;
		12'd0658: rd_data_0 <= 24'h7e007f;
		12'd0659: rd_data_0 <= 24'h7e007f;
		12'd0660: rd_data_0 <= 24'h7f007f;
		12'd0661: rd_data_0 <= 24'h7f007f;
		12'd0662: rd_data_0 <= 24'h7f007f;
		12'd0663: rd_data_0 <= 24'h7f007f;
		12'd0664: rd_data_0 <= 24'h7f007f;
		12'd0665: rd_data_0 <= 24'h7f007f;
		12'd0666: rd_data_0 <= 24'h7f007f;
		12'd0667: rd_data_0 <= 24'h7f007f;
		12'd0668: rd_data_0 <= 24'h7f007f;
		12'd0669: rd_data_0 <= 24'h7f007f;
		12'd0670: rd_data_0 <= 24'h7f007f;
		12'd0671: rd_data_0 <= 24'h7f007f;
		12'd0672: rd_data_0 <= 24'h7f007f;
		12'd0673: rd_data_0 <= 24'h7f007f;
		12'd0674: rd_data_0 <= 24'h7f007f;
		12'd0675: rd_data_0 <= 24'h7f007f;
		12'd0676: rd_data_0 <= 24'h7f007f;
		12'd0677: rd_data_0 <= 24'h7f007f;
		12'd0678: rd_data_0 <= 24'h7f007f;
		12'd0679: rd_data_0 <= 24'h7f007f;
		12'd0680: rd_data_0 <= 24'h7f007f;
		12'd0681: rd_data_0 <= 24'h7f007f;
		12'd0682: rd_data_0 <= 24'h7f007f;
		12'd0683: rd_data_0 <= 24'h7f007f;
		12'd0684: rd_data_0 <= 24'h7f007f;
		12'd0685: rd_data_0 <= 24'h7f007f;
		12'd0686: rd_data_0 <= 24'h7f007f;
		12'd0687: rd_data_0 <= 24'h7f007f;
		12'd0688: rd_data_0 <= 24'h7f007f;
		12'd0689: rd_data_0 <= 24'h7f007f;
		12'd0690: rd_data_0 <= 24'h7f007f;
		12'd0691: rd_data_0 <= 24'h7f007f;
		12'd0692: rd_data_0 <= 24'h7f007f;
		12'd0693: rd_data_0 <= 24'h7f007f;
		12'd0694: rd_data_0 <= 24'h7f007f;
		12'd0695: rd_data_0 <= 24'h7f007f;
		12'd0696: rd_data_0 <= 24'h7f007f;
		12'd0697: rd_data_0 <= 24'h7f007f;
		12'd0698: rd_data_0 <= 24'h7f007f;
		12'd0699: rd_data_0 <= 24'h7f007f;
		12'd0700: rd_data_0 <= 24'h7f007f;
		12'd0701: rd_data_0 <= 24'h7f007f;
		12'd0702: rd_data_0 <= 24'h7f007f;
		12'd0703: rd_data_0 <= 24'h7f007f;
		12'd0704: rd_data_0 <= 24'h81007d;
		12'd0705: rd_data_0 <= 24'h81007d;
		12'd0706: rd_data_0 <= 24'h81007d;
		12'd0707: rd_data_0 <= 24'h81007d;
		12'd0708: rd_data_0 <= 24'h81007f;
		12'd0709: rd_data_0 <= 24'h81007f;
		12'd0710: rd_data_0 <= 24'h7f007f;
		12'd0711: rd_data_0 <= 24'h7f007f;
		12'd0712: rd_data_0 <= 24'h7e007f;
		12'd0713: rd_data_0 <= 24'h7e007f;
		12'd0714: rd_data_0 <= 24'h7c017f;
		12'd0715: rd_data_0 <= 24'h7c017f;
		12'd0716: rd_data_0 <= 24'h7e007f;
		12'd0717: rd_data_0 <= 24'h7e007f;
		12'd0718: rd_data_0 <= 24'h7e007f;
		12'd0719: rd_data_0 <= 24'h7e007f;
		12'd0720: rd_data_0 <= 24'h7e007f;
		12'd0721: rd_data_0 <= 24'h7e007f;
		12'd0722: rd_data_0 <= 24'h7e007f;
		12'd0723: rd_data_0 <= 24'h7e007f;
		12'd0724: rd_data_0 <= 24'h7f007f;
		12'd0725: rd_data_0 <= 24'h7f007f;
		12'd0726: rd_data_0 <= 24'h7f007f;
		12'd0727: rd_data_0 <= 24'h7f007f;
		12'd0728: rd_data_0 <= 24'h7f007f;
		12'd0729: rd_data_0 <= 24'h7f007f;
		12'd0730: rd_data_0 <= 24'h7f007f;
		12'd0731: rd_data_0 <= 24'h7f007f;
		12'd0732: rd_data_0 <= 24'h7f007f;
		12'd0733: rd_data_0 <= 24'h7f007f;
		12'd0734: rd_data_0 <= 24'h7f007f;
		12'd0735: rd_data_0 <= 24'h7f007f;
		12'd0736: rd_data_0 <= 24'h7f007f;
		12'd0737: rd_data_0 <= 24'h7f007f;
		12'd0738: rd_data_0 <= 24'h7f007f;
		12'd0739: rd_data_0 <= 24'h7f007f;
		12'd0740: rd_data_0 <= 24'h7f007f;
		12'd0741: rd_data_0 <= 24'h7f007f;
		12'd0742: rd_data_0 <= 24'h7f007f;
		12'd0743: rd_data_0 <= 24'h7f007f;
		12'd0744: rd_data_0 <= 24'h7f007f;
		12'd0745: rd_data_0 <= 24'h7f007f;
		12'd0746: rd_data_0 <= 24'h7f007f;
		12'd0747: rd_data_0 <= 24'h7f007f;
		12'd0748: rd_data_0 <= 24'h7f007f;
		12'd0749: rd_data_0 <= 24'h7f007f;
		12'd0750: rd_data_0 <= 24'h7f007f;
		12'd0751: rd_data_0 <= 24'h7f007f;
		12'd0752: rd_data_0 <= 24'h7f007f;
		12'd0753: rd_data_0 <= 24'h7f007f;
		12'd0754: rd_data_0 <= 24'h7f007f;
		12'd0755: rd_data_0 <= 24'h7f007f;
		12'd0756: rd_data_0 <= 24'h7f007f;
		12'd0757: rd_data_0 <= 24'h7f007f;
		12'd0758: rd_data_0 <= 24'h7f007f;
		12'd0759: rd_data_0 <= 24'h7f007f;
		12'd0760: rd_data_0 <= 24'h7f007f;
		12'd0761: rd_data_0 <= 24'h7f007f;
		12'd0762: rd_data_0 <= 24'h7f007f;
		12'd0763: rd_data_0 <= 24'h7f007f;
		12'd0764: rd_data_0 <= 24'h7f007f;
		12'd0765: rd_data_0 <= 24'h7f007f;
		12'd0766: rd_data_0 <= 24'h7f007f;
		12'd0767: rd_data_0 <= 24'h7f007f;
		12'd0768: rd_data_0 <= 24'h81007d;
		12'd0769: rd_data_0 <= 24'h81007d;
		12'd0770: rd_data_0 <= 24'h81007d;
		12'd0771: rd_data_0 <= 24'h81007d;
		12'd0772: rd_data_0 <= 24'h81007f;
		12'd0773: rd_data_0 <= 24'h81007f;
		12'd0774: rd_data_0 <= 24'h7f007f;
		12'd0775: rd_data_0 <= 24'h7f007f;
		12'd0776: rd_data_0 <= 24'h7e007f;
		12'd0777: rd_data_0 <= 24'h7e007f;
		12'd0778: rd_data_0 <= 24'h7e007f;
		12'd0779: rd_data_0 <= 24'h7e007f;
		12'd0780: rd_data_0 <= 24'h7e0081;
		12'd0781: rd_data_0 <= 24'h7e0081;
		12'd0782: rd_data_0 <= 24'h7e0081;
		12'd0783: rd_data_0 <= 24'h7e0081;
		12'd0784: rd_data_0 <= 24'h7e007f;
		12'd0785: rd_data_0 <= 24'h7e007f;
		12'd0786: rd_data_0 <= 24'h7e007f;
		12'd0787: rd_data_0 <= 24'h7e007f;
		12'd0788: rd_data_0 <= 24'h7f007f;
		12'd0789: rd_data_0 <= 24'h7f007f;
		12'd0790: rd_data_0 <= 24'h7f007f;
		12'd0791: rd_data_0 <= 24'h7f007f;
		12'd0792: rd_data_0 <= 24'h7f007f;
		12'd0793: rd_data_0 <= 24'h7f007f;
		12'd0794: rd_data_0 <= 24'h7f007f;
		12'd0795: rd_data_0 <= 24'h7f007f;
		12'd0796: rd_data_0 <= 24'h7f007f;
		12'd0797: rd_data_0 <= 24'h7f007f;
		12'd0798: rd_data_0 <= 24'h7f007f;
		12'd0799: rd_data_0 <= 24'h7f007f;
		12'd0800: rd_data_0 <= 24'h7f007f;
		12'd0801: rd_data_0 <= 24'h7f007f;
		12'd0802: rd_data_0 <= 24'h7f007f;
		12'd0803: rd_data_0 <= 24'h7f007f;
		12'd0804: rd_data_0 <= 24'h7f007f;
		12'd0805: rd_data_0 <= 24'h7f007f;
		12'd0806: rd_data_0 <= 24'h7f007f;
		12'd0807: rd_data_0 <= 24'h7f007f;
		12'd0808: rd_data_0 <= 24'h7f007f;
		12'd0809: rd_data_0 <= 24'h7f007f;
		12'd0810: rd_data_0 <= 24'h7f007f;
		12'd0811: rd_data_0 <= 24'h7f007f;
		12'd0812: rd_data_0 <= 24'h7f007f;
		12'd0813: rd_data_0 <= 24'h7f007f;
		12'd0814: rd_data_0 <= 24'h7f007f;
		12'd0815: rd_data_0 <= 24'h7f007f;
		12'd0816: rd_data_0 <= 24'h7f007f;
		12'd0817: rd_data_0 <= 24'h7f007f;
		12'd0818: rd_data_0 <= 24'h7f007f;
		12'd0819: rd_data_0 <= 24'h7f007f;
		12'd0820: rd_data_0 <= 24'h7f007f;
		12'd0821: rd_data_0 <= 24'h7f007f;
		12'd0822: rd_data_0 <= 24'h7f007f;
		12'd0823: rd_data_0 <= 24'h7f007f;
		12'd0824: rd_data_0 <= 24'h7f007f;
		12'd0825: rd_data_0 <= 24'h7f007f;
		12'd0826: rd_data_0 <= 24'h7f007f;
		12'd0827: rd_data_0 <= 24'h7f007f;
		12'd0828: rd_data_0 <= 24'h7f007f;
		12'd0829: rd_data_0 <= 24'h7f007f;
		12'd0830: rd_data_0 <= 24'h7f007f;
		12'd0831: rd_data_0 <= 24'h7f007f;
		12'd0832: rd_data_0 <= 24'h81007d;
		12'd0833: rd_data_0 <= 24'h81007d;
		12'd0834: rd_data_0 <= 24'h81007d;
		12'd0835: rd_data_0 <= 24'h81007d;
		12'd0836: rd_data_0 <= 24'h81007f;
		12'd0837: rd_data_0 <= 24'h81007f;
		12'd0838: rd_data_0 <= 24'h7f007f;
		12'd0839: rd_data_0 <= 24'h7f007f;
		12'd0840: rd_data_0 <= 24'h7e007f;
		12'd0841: rd_data_0 <= 24'h7e007f;
		12'd0842: rd_data_0 <= 24'h7e007f;
		12'd0843: rd_data_0 <= 24'h7e007f;
		12'd0844: rd_data_0 <= 24'h7e0081;
		12'd0845: rd_data_0 <= 24'h7e0081;
		12'd0846: rd_data_0 <= 24'h7e0081;
		12'd0847: rd_data_0 <= 24'h7e0081;
		12'd0848: rd_data_0 <= 24'h7e007f;
		12'd0849: rd_data_0 <= 24'h7e007f;
		12'd0850: rd_data_0 <= 24'h7e007f;
		12'd0851: rd_data_0 <= 24'h7e007f;
		12'd0852: rd_data_0 <= 24'h7f007f;
		12'd0853: rd_data_0 <= 24'h7f007f;
		12'd0854: rd_data_0 <= 24'h7f007f;
		12'd0855: rd_data_0 <= 24'h7f007f;
		12'd0856: rd_data_0 <= 24'h7f007f;
		12'd0857: rd_data_0 <= 24'h7f007f;
		12'd0858: rd_data_0 <= 24'h7f007f;
		12'd0859: rd_data_0 <= 24'h7f007f;
		12'd0860: rd_data_0 <= 24'h7f007f;
		12'd0861: rd_data_0 <= 24'h7f007f;
		12'd0862: rd_data_0 <= 24'h7f007f;
		12'd0863: rd_data_0 <= 24'h7f007f;
		12'd0864: rd_data_0 <= 24'h7f007f;
		12'd0865: rd_data_0 <= 24'h7f007f;
		12'd0866: rd_data_0 <= 24'h7f007f;
		12'd0867: rd_data_0 <= 24'h7f007f;
		12'd0868: rd_data_0 <= 24'h7f007f;
		12'd0869: rd_data_0 <= 24'h7f007f;
		12'd0870: rd_data_0 <= 24'h7f007f;
		12'd0871: rd_data_0 <= 24'h7f007f;
		12'd0872: rd_data_0 <= 24'h7f007f;
		12'd0873: rd_data_0 <= 24'h7f007f;
		12'd0874: rd_data_0 <= 24'h7f007f;
		12'd0875: rd_data_0 <= 24'h7f007f;
		12'd0876: rd_data_0 <= 24'h7f007f;
		12'd0877: rd_data_0 <= 24'h7f007f;
		12'd0878: rd_data_0 <= 24'h7f007f;
		12'd0879: rd_data_0 <= 24'h7f007f;
		12'd0880: rd_data_0 <= 24'h7f007f;
		12'd0881: rd_data_0 <= 24'h7f007f;
		12'd0882: rd_data_0 <= 24'h7f007f;
		12'd0883: rd_data_0 <= 24'h7f007f;
		12'd0884: rd_data_0 <= 24'h7f007f;
		12'd0885: rd_data_0 <= 24'h7f007f;
		12'd0886: rd_data_0 <= 24'h7f007f;
		12'd0887: rd_data_0 <= 24'h7f007f;
		12'd0888: rd_data_0 <= 24'h7f007f;
		12'd0889: rd_data_0 <= 24'h7f007f;
		12'd0890: rd_data_0 <= 24'h7f007f;
		12'd0891: rd_data_0 <= 24'h7f007f;
		12'd0892: rd_data_0 <= 24'h7f007f;
		12'd0893: rd_data_0 <= 24'h7f007f;
		12'd0894: rd_data_0 <= 24'h7f007f;
		12'd0895: rd_data_0 <= 24'h7f007f;
		12'd0896: rd_data_0 <= 24'h81007d;
		12'd0897: rd_data_0 <= 24'h81007d;
		12'd0898: rd_data_0 <= 24'h81007d;
		12'd0899: rd_data_0 <= 24'h81007d;
		12'd0900: rd_data_0 <= 24'h81007f;
		12'd0901: rd_data_0 <= 24'h81007f;
		12'd0902: rd_data_0 <= 24'h7f007f;
		12'd0903: rd_data_0 <= 24'h7f007f;
		12'd0904: rd_data_0 <= 24'h7e007f;
		12'd0905: rd_data_0 <= 24'h7e007f;
		12'd0906: rd_data_0 <= 24'h7e007f;
		12'd0907: rd_data_0 <= 24'h7e007f;
		12'd0908: rd_data_0 <= 24'h7e0081;
		12'd0909: rd_data_0 <= 24'h7e0081;
		12'd0910: rd_data_0 <= 24'h7e0081;
		12'd0911: rd_data_0 <= 24'h7e0081;
		12'd0912: rd_data_0 <= 24'h7e007f;
		12'd0913: rd_data_0 <= 24'h7e007f;
		12'd0914: rd_data_0 <= 24'h7e007f;
		12'd0915: rd_data_0 <= 24'h7e007f;
		12'd0916: rd_data_0 <= 24'h7f007f;
		12'd0917: rd_data_0 <= 24'h7f007f;
		12'd0918: rd_data_0 <= 24'h7f007f;
		12'd0919: rd_data_0 <= 24'h7f007f;
		12'd0920: rd_data_0 <= 24'h7f007f;
		12'd0921: rd_data_0 <= 24'h7f007f;
		12'd0922: rd_data_0 <= 24'h7f007f;
		12'd0923: rd_data_0 <= 24'h7f007f;
		12'd0924: rd_data_0 <= 24'h7f007f;
		12'd0925: rd_data_0 <= 24'h7f007f;
		12'd0926: rd_data_0 <= 24'h7f007f;
		12'd0927: rd_data_0 <= 24'h7f007f;
		12'd0928: rd_data_0 <= 24'h7f007f;
		12'd0929: rd_data_0 <= 24'h7f007f;
		12'd0930: rd_data_0 <= 24'h7f007f;
		12'd0931: rd_data_0 <= 24'h7f007f;
		12'd0932: rd_data_0 <= 24'h7f007f;
		12'd0933: rd_data_0 <= 24'h7f007f;
		12'd0934: rd_data_0 <= 24'h7f007f;
		12'd0935: rd_data_0 <= 24'h7f007f;
		12'd0936: rd_data_0 <= 24'h7f0080;
		12'd0937: rd_data_0 <= 24'h7f0080;
		12'd0938: rd_data_0 <= 24'h7f007f;
		12'd0939: rd_data_0 <= 24'h7f007f;
		12'd0940: rd_data_0 <= 24'h7f007f;
		12'd0941: rd_data_0 <= 24'h7f007f;
		12'd0942: rd_data_0 <= 24'h7f007f;
		12'd0943: rd_data_0 <= 24'h7e007f;
		12'd0944: rd_data_0 <= 24'h7e007f;
		12'd0945: rd_data_0 <= 24'h7f007f;
		12'd0946: rd_data_0 <= 24'h7f007f;
		12'd0947: rd_data_0 <= 24'h7f007f;
		12'd0948: rd_data_0 <= 24'h7f007f;
		12'd0949: rd_data_0 <= 24'h7f007f;
		12'd0950: rd_data_0 <= 24'h7f007f;
		12'd0951: rd_data_0 <= 24'h7f007f;
		12'd0952: rd_data_0 <= 24'h7f007f;
		12'd0953: rd_data_0 <= 24'h7f007f;
		12'd0954: rd_data_0 <= 24'h7f007f;
		12'd0955: rd_data_0 <= 24'h7f007f;
		12'd0956: rd_data_0 <= 24'h7f007f;
		12'd0957: rd_data_0 <= 24'h7f007f;
		12'd0958: rd_data_0 <= 24'h7f007f;
		12'd0959: rd_data_0 <= 24'h7f007f;
		12'd0960: rd_data_0 <= 24'h81007d;
		12'd0961: rd_data_0 <= 24'h81007d;
		12'd0962: rd_data_0 <= 24'h81007d;
		12'd0963: rd_data_0 <= 24'h81007d;
		12'd0964: rd_data_0 <= 24'h81007f;
		12'd0965: rd_data_0 <= 24'h81007f;
		12'd0966: rd_data_0 <= 24'h7f007f;
		12'd0967: rd_data_0 <= 24'h7f007f;
		12'd0968: rd_data_0 <= 24'h7e007f;
		12'd0969: rd_data_0 <= 24'h7e007f;
		12'd0970: rd_data_0 <= 24'h7e007f;
		12'd0971: rd_data_0 <= 24'h7e007f;
		12'd0972: rd_data_0 <= 24'h7e0081;
		12'd0973: rd_data_0 <= 24'h7e0081;
		12'd0974: rd_data_0 <= 24'h7e0081;
		12'd0975: rd_data_0 <= 24'h7e0081;
		12'd0976: rd_data_0 <= 24'h7d017f;
		12'd0977: rd_data_0 <= 24'h7d017f;
		12'd0978: rd_data_0 <= 24'h7e007f;
		12'd0979: rd_data_0 <= 24'h7e007f;
		12'd0980: rd_data_0 <= 24'h7e007f;
		12'd0981: rd_data_0 <= 24'h7e007f;
		12'd0982: rd_data_0 <= 24'h80007f;
		12'd0983: rd_data_0 <= 24'h82007f;
		12'd0984: rd_data_0 <= 24'h81007f;
		12'd0985: rd_data_0 <= 24'h800080;
		12'd0986: rd_data_0 <= 24'h800080;
		12'd0987: rd_data_0 <= 24'h80007e;
		12'd0988: rd_data_0 <= 24'h7e007d;
		12'd0989: rd_data_0 <= 24'h7e007e;
		12'd0990: rd_data_0 <= 24'h800180;
		12'd0991: rd_data_0 <= 24'h820181;
		12'd0992: rd_data_0 <= 24'h800080;
		12'd0993: rd_data_0 <= 24'h7e007f;
		12'd0994: rd_data_0 <= 24'h7e007f;
		12'd0995: rd_data_0 <= 24'h7e007e;
		12'd0996: rd_data_0 <= 24'h7e017e;
		12'd0997: rd_data_0 <= 24'h7f017d;
		12'd0998: rd_data_0 <= 24'h7e017c;
		12'd0999: rd_data_0 <= 24'h7d007c;
		12'd1000: rd_data_0 <= 24'h7c027a;
		12'd1001: rd_data_0 <= 24'h7b0378;
		12'd1002: rd_data_0 <= 24'h7d027b;
		12'd1003: rd_data_0 <= 24'h80007d;
		12'd1004: rd_data_0 <= 24'h810080;
		12'd1005: rd_data_0 <= 24'h7f0080;
		12'd1006: rd_data_0 <= 24'h7e0080;
		12'd1007: rd_data_0 <= 24'h7c017f;
		12'd1008: rd_data_0 <= 24'h7c017f;
		12'd1009: rd_data_0 <= 24'h7e007f;
		12'd1010: rd_data_0 <= 24'h7f007f;
		12'd1011: rd_data_0 <= 24'h7f007f;
		12'd1012: rd_data_0 <= 24'h7f007f;
		12'd1013: rd_data_0 <= 24'h7f007f;
		12'd1014: rd_data_0 <= 24'h7f007f;
		12'd1015: rd_data_0 <= 24'h7f007f;
		12'd1016: rd_data_0 <= 24'h7f007f;
		12'd1017: rd_data_0 <= 24'h7f007f;
		12'd1018: rd_data_0 <= 24'h7f007f;
		12'd1019: rd_data_0 <= 24'h7f007f;
		12'd1020: rd_data_0 <= 24'h7f007f;
		12'd1021: rd_data_0 <= 24'h7f007f;
		12'd1022: rd_data_0 <= 24'h7f007f;
		12'd1023: rd_data_0 <= 24'h7f007f;
		12'd1024: rd_data_0 <= 24'h7f007f;
		12'd1025: rd_data_0 <= 24'h7f007f;
		12'd1026: rd_data_0 <= 24'h7f007f;
		12'd1027: rd_data_0 <= 24'h7f007f;
		12'd1028: rd_data_0 <= 24'h7f007f;
		12'd1029: rd_data_0 <= 24'h7f007f;
		12'd1030: rd_data_0 <= 24'h7f007f;
		12'd1031: rd_data_0 <= 24'h7f007f;
		12'd1032: rd_data_0 <= 24'h7f007f;
		12'd1033: rd_data_0 <= 24'h7f007f;
		12'd1034: rd_data_0 <= 24'h7e007f;
		12'd1035: rd_data_0 <= 24'h7e007f;
		12'd1036: rd_data_0 <= 24'h7f007f;
		12'd1037: rd_data_0 <= 24'h7f007f;
		12'd1038: rd_data_0 <= 24'h7f007f;
		12'd1039: rd_data_0 <= 24'h7d017f;
		12'd1040: rd_data_0 <= 24'h79037f;
		12'd1041: rd_data_0 <= 24'h79047d;
		12'd1042: rd_data_0 <= 24'h80017d;
		12'd1043: rd_data_0 <= 24'h83007d;
		12'd1044: rd_data_0 <= 24'h7e017d;
		12'd1045: rd_data_0 <= 24'h7c027d;
		12'd1046: rd_data_0 <= 24'h81017d;
		12'd1047: rd_data_0 <= 24'h86007f;
		12'd1048: rd_data_0 <= 24'h860084;
		12'd1049: rd_data_0 <= 24'h840085;
		12'd1050: rd_data_0 <= 24'h830081;
		12'd1051: rd_data_0 <= 24'h80007c;
		12'd1052: rd_data_0 <= 24'h81057e;
		12'd1053: rd_data_0 <= 24'h7c047b;
		12'd1054: rd_data_0 <= 24'h80007f;
		12'd1055: rd_data_0 <= 24'h8b0088;
		12'd1056: rd_data_0 <= 24'h8a038a;
		12'd1057: rd_data_0 <= 24'h850689;
		12'd1058: rd_data_0 <= 24'h800283;
		12'd1059: rd_data_0 <= 24'h7e017d;
		12'd1060: rd_data_0 <= 24'h7c0078;
		12'd1061: rd_data_0 <= 24'h7a0074;
		12'd1062: rd_data_0 <= 24'h7e0275;
		12'd1063: rd_data_0 <= 24'h7d0472;
		12'd1064: rd_data_0 <= 24'h76076c;
		12'd1065: rd_data_0 <= 24'h730e6b;
		12'd1066: rd_data_0 <= 24'h74036b;
		12'd1067: rd_data_0 <= 24'h810077;
		12'd1068: rd_data_0 <= 24'h80007e;
		12'd1069: rd_data_0 <= 24'h7e0086;
		12'd1070: rd_data_0 <= 24'h7c0184;
		12'd1071: rd_data_0 <= 24'h7b0280;
		12'd1072: rd_data_0 <= 24'h7c017f;
		12'd1073: rd_data_0 <= 24'h7e007f;
		12'd1074: rd_data_0 <= 24'h7f007f;
		12'd1075: rd_data_0 <= 24'h7f007f;
		12'd1076: rd_data_0 <= 24'h7f007f;
		12'd1077: rd_data_0 <= 24'h7f007f;
		12'd1078: rd_data_0 <= 24'h7f007f;
		12'd1079: rd_data_0 <= 24'h7f007f;
		12'd1080: rd_data_0 <= 24'h7f007f;
		12'd1081: rd_data_0 <= 24'h7f007f;
		12'd1082: rd_data_0 <= 24'h7f007f;
		12'd1083: rd_data_0 <= 24'h7f007f;
		12'd1084: rd_data_0 <= 24'h7f007f;
		12'd1085: rd_data_0 <= 24'h7f007f;
		12'd1086: rd_data_0 <= 24'h7f007f;
		12'd1087: rd_data_0 <= 24'h7f007f;
		12'd1088: rd_data_0 <= 24'h7f007f;
		12'd1089: rd_data_0 <= 24'h7f007f;
		12'd1090: rd_data_0 <= 24'h7f007f;
		12'd1091: rd_data_0 <= 24'h7f007f;
		12'd1092: rd_data_0 <= 24'h7f007f;
		12'd1093: rd_data_0 <= 24'h7f007f;
		12'd1094: rd_data_0 <= 24'h7f007f;
		12'd1095: rd_data_0 <= 24'h7f007f;
		12'd1096: rd_data_0 <= 24'h7f007f;
		12'd1097: rd_data_0 <= 24'h7f007f;
		12'd1098: rd_data_0 <= 24'h7e007f;
		12'd1099: rd_data_0 <= 24'h7e007f;
		12'd1100: rd_data_0 <= 24'h7f007f;
		12'd1101: rd_data_0 <= 24'h7f007f;
		12'd1102: rd_data_0 <= 24'h7f007f;
		12'd1103: rd_data_0 <= 24'h7f007f;
		12'd1104: rd_data_0 <= 24'h79027f;
		12'd1105: rd_data_0 <= 24'h79037e;
		12'd1106: rd_data_0 <= 24'h82007e;
		12'd1107: rd_data_0 <= 24'h85007e;
		12'd1108: rd_data_0 <= 24'h7e017e;
		12'd1109: rd_data_0 <= 24'h7a027e;
		12'd1110: rd_data_0 <= 24'h81017e;
		12'd1111: rd_data_0 <= 24'h860080;
		12'd1112: rd_data_0 <= 24'h870086;
		12'd1113: rd_data_0 <= 24'h850088;
		12'd1114: rd_data_0 <= 24'h840083;
		12'd1115: rd_data_0 <= 24'h7f007d;
		12'd1116: rd_data_0 <= 24'h790177;
		12'd1117: rd_data_0 <= 24'h750173;
		12'd1118: rd_data_0 <= 24'h7f017e;
		12'd1119: rd_data_0 <= 24'h850085;
		12'd1120: rd_data_0 <= 24'h7e0381;
		12'd1121: rd_data_0 <= 24'h710479;
		12'd1122: rd_data_0 <= 24'h68006f;
		12'd1123: rd_data_0 <= 24'h710974;
		12'd1124: rd_data_0 <= 24'h730d72;
		12'd1125: rd_data_0 <= 24'h710b6a;
		12'd1126: rd_data_0 <= 24'h79136f;
		12'd1127: rd_data_0 <= 24'h700f65;
		12'd1128: rd_data_0 <= 24'h621356;
		12'd1129: rd_data_0 <= 24'h602356;
		12'd1130: rd_data_0 <= 24'h6b2062;
		12'd1131: rd_data_0 <= 24'h710969;
		12'd1132: rd_data_0 <= 24'h710070;
		12'd1133: rd_data_0 <= 24'h780381;
		12'd1134: rd_data_0 <= 24'h790381;
		12'd1135: rd_data_0 <= 24'h7b037e;
		12'd1136: rd_data_0 <= 24'h7c027e;
		12'd1137: rd_data_0 <= 24'h7e007f;
		12'd1138: rd_data_0 <= 24'h7f007f;
		12'd1139: rd_data_0 <= 24'h7f007f;
		12'd1140: rd_data_0 <= 24'h7f007f;
		12'd1141: rd_data_0 <= 24'h7f007f;
		12'd1142: rd_data_0 <= 24'h7f007f;
		12'd1143: rd_data_0 <= 24'h7f007f;
		12'd1144: rd_data_0 <= 24'h7f007f;
		12'd1145: rd_data_0 <= 24'h7f007f;
		12'd1146: rd_data_0 <= 24'h7f007f;
		12'd1147: rd_data_0 <= 24'h7f007f;
		12'd1148: rd_data_0 <= 24'h7f007f;
		12'd1149: rd_data_0 <= 24'h7f007f;
		12'd1150: rd_data_0 <= 24'h7f007f;
		12'd1151: rd_data_0 <= 24'h7f007f;
		12'd1152: rd_data_0 <= 24'h7f007f;
		12'd1153: rd_data_0 <= 24'h7f007f;
		12'd1154: rd_data_0 <= 24'h7f007f;
		12'd1155: rd_data_0 <= 24'h7f007f;
		12'd1156: rd_data_0 <= 24'h7f007f;
		12'd1157: rd_data_0 <= 24'h7f007f;
		12'd1158: rd_data_0 <= 24'h7f007f;
		12'd1159: rd_data_0 <= 24'h7f007f;
		12'd1160: rd_data_0 <= 24'h7f007f;
		12'd1161: rd_data_0 <= 24'h7f007f;
		12'd1162: rd_data_0 <= 24'h7e0081;
		12'd1163: rd_data_0 <= 24'h7e0081;
		12'd1164: rd_data_0 <= 24'h7f0081;
		12'd1165: rd_data_0 <= 24'h7f0081;
		12'd1166: rd_data_0 <= 24'h7f0081;
		12'd1167: rd_data_0 <= 24'h7f0081;
		12'd1168: rd_data_0 <= 24'h7d0081;
		12'd1169: rd_data_0 <= 24'h7d0081;
		12'd1170: rd_data_0 <= 24'h830082;
		12'd1171: rd_data_0 <= 24'h850082;
		12'd1172: rd_data_0 <= 24'h7d0082;
		12'd1173: rd_data_0 <= 24'h790383;
		12'd1174: rd_data_0 <= 24'h7c0184;
		12'd1175: rd_data_0 <= 24'h800084;
		12'd1176: rd_data_0 <= 24'h830085;
		12'd1177: rd_data_0 <= 24'h830086;
		12'd1178: rd_data_0 <= 24'h7f0086;
		12'd1179: rd_data_0 <= 24'h7e0185;
		12'd1180: rd_data_0 <= 24'h800284;
		12'd1181: rd_data_0 <= 24'h800380;
		12'd1182: rd_data_0 <= 24'h770379;
		12'd1183: rd_data_0 <= 24'h6b0571;
		12'd1184: rd_data_0 <= 24'h62116e;
		12'd1185: rd_data_0 <= 24'h541564;
		12'd1186: rd_data_0 <= 24'h4a1259;
		12'd1187: rd_data_0 <= 24'h50195b;
		12'd1188: rd_data_0 <= 24'h511a57;
		12'd1189: rd_data_0 <= 24'h501a51;
		12'd1190: rd_data_0 <= 24'h551f52;
		12'd1191: rd_data_0 <= 24'h52224e;
		12'd1192: rd_data_0 <= 24'h4d3748;
		12'd1193: rd_data_0 <= 24'h5b6055;
		12'd1194: rd_data_0 <= 24'h6f6a6d;
		12'd1195: rd_data_0 <= 24'h1c001d;
		12'd1196: rd_data_0 <= 24'h410041;
		12'd1197: rd_data_0 <= 24'h6e0d6c;
		12'd1198: rd_data_0 <= 24'h780776;
		12'd1199: rd_data_0 <= 24'h7a0478;
		12'd1200: rd_data_0 <= 24'h7d027a;
		12'd1201: rd_data_0 <= 24'h7e017e;
		12'd1202: rd_data_0 <= 24'h7f007f;
		12'd1203: rd_data_0 <= 24'h7f007f;
		12'd1204: rd_data_0 <= 24'h7f007f;
		12'd1205: rd_data_0 <= 24'h7f007f;
		12'd1206: rd_data_0 <= 24'h7f007f;
		12'd1207: rd_data_0 <= 24'h7f007f;
		12'd1208: rd_data_0 <= 24'h7f007f;
		12'd1209: rd_data_0 <= 24'h7f007f;
		12'd1210: rd_data_0 <= 24'h7f007f;
		12'd1211: rd_data_0 <= 24'h7f007f;
		12'd1212: rd_data_0 <= 24'h7f007f;
		12'd1213: rd_data_0 <= 24'h7f007f;
		12'd1214: rd_data_0 <= 24'h7f007f;
		12'd1215: rd_data_0 <= 24'h7f007f;
		12'd1216: rd_data_0 <= 24'h7f007f;
		12'd1217: rd_data_0 <= 24'h7f007f;
		12'd1218: rd_data_0 <= 24'h7f007f;
		12'd1219: rd_data_0 <= 24'h7f007f;
		12'd1220: rd_data_0 <= 24'h7f007f;
		12'd1221: rd_data_0 <= 24'h7f007f;
		12'd1222: rd_data_0 <= 24'h7f007f;
		12'd1223: rd_data_0 <= 24'h7f007f;
		12'd1224: rd_data_0 <= 24'h7f007f;
		12'd1225: rd_data_0 <= 24'h7f007f;
		12'd1226: rd_data_0 <= 24'h7e0081;
		12'd1227: rd_data_0 <= 24'h7e0081;
		12'd1228: rd_data_0 <= 24'h7f0081;
		12'd1229: rd_data_0 <= 24'h7f0081;
		12'd1230: rd_data_0 <= 24'h7f0081;
		12'd1231: rd_data_0 <= 24'h7f0081;
		12'd1232: rd_data_0 <= 24'h7f0082;
		12'd1233: rd_data_0 <= 24'h7f0081;
		12'd1234: rd_data_0 <= 24'h810084;
		12'd1235: rd_data_0 <= 24'h820083;
		12'd1236: rd_data_0 <= 24'h7b0082;
		12'd1237: rd_data_0 <= 24'h790284;
		12'd1238: rd_data_0 <= 24'h7b0286;
		12'd1239: rd_data_0 <= 24'h7c0185;
		12'd1240: rd_data_0 <= 24'h7e0083;
		12'd1241: rd_data_0 <= 24'h7f0082;
		12'd1242: rd_data_0 <= 24'h7d0083;
		12'd1243: rd_data_0 <= 24'h790284;
		12'd1244: rd_data_0 <= 24'h7b0782;
		12'd1245: rd_data_0 <= 24'h730773;
		12'd1246: rd_data_0 <= 24'h5c0960;
		12'd1247: rd_data_0 <= 24'h622c6a;
		12'd1248: rd_data_0 <= 24'h6d507b;
		12'd1249: rd_data_0 <= 24'h695d7c;
		12'd1250: rd_data_0 <= 24'h655c75;
		12'd1251: rd_data_0 <= 24'h50485c;
		12'd1252: rd_data_0 <= 24'h3f3846;
		12'd1253: rd_data_0 <= 24'h423c44;
		12'd1254: rd_data_0 <= 24'h40393f;
		12'd1255: rd_data_0 <= 24'h5b5c59;
		12'd1256: rd_data_0 <= 24'h738c6f;
		12'd1257: rd_data_0 <= 24'h50824c;
		12'd1258: rd_data_0 <= 24'h507d52;
		12'd1259: rd_data_0 <= 24'h36463d;
		12'd1260: rd_data_0 <= 24'h5d3d5e;
		12'd1261: rd_data_0 <= 24'h580851;
		12'd1262: rd_data_0 <= 24'h73086b;
		12'd1263: rd_data_0 <= 24'h780375;
		12'd1264: rd_data_0 <= 24'h7d027c;
		12'd1265: rd_data_0 <= 24'h7e007f;
		12'd1266: rd_data_0 <= 24'h7f007f;
		12'd1267: rd_data_0 <= 24'h7f007f;
		12'd1268: rd_data_0 <= 24'h7f007f;
		12'd1269: rd_data_0 <= 24'h7f007f;
		12'd1270: rd_data_0 <= 24'h7f007f;
		12'd1271: rd_data_0 <= 24'h7f007f;
		12'd1272: rd_data_0 <= 24'h7f007f;
		12'd1273: rd_data_0 <= 24'h7f007f;
		12'd1274: rd_data_0 <= 24'h7f007f;
		12'd1275: rd_data_0 <= 24'h7f007f;
		12'd1276: rd_data_0 <= 24'h7f007f;
		12'd1277: rd_data_0 <= 24'h7f007f;
		12'd1278: rd_data_0 <= 24'h7f007f;
		12'd1279: rd_data_0 <= 24'h7f007f;
		12'd1280: rd_data_0 <= 24'h7f007f;
		12'd1281: rd_data_0 <= 24'h7f007f;
		12'd1282: rd_data_0 <= 24'h7f007f;
		12'd1283: rd_data_0 <= 24'h7f007f;
		12'd1284: rd_data_0 <= 24'h7f007f;
		12'd1285: rd_data_0 <= 24'h7f007f;
		12'd1286: rd_data_0 <= 24'h7f007f;
		12'd1287: rd_data_0 <= 24'h7f007f;
		12'd1288: rd_data_0 <= 24'h7f007f;
		12'd1289: rd_data_0 <= 24'h7f007f;
		12'd1290: rd_data_0 <= 24'h7f0080;
		12'd1291: rd_data_0 <= 24'h7f0080;
		12'd1292: rd_data_0 <= 24'h7f0080;
		12'd1293: rd_data_0 <= 24'h7f0080;
		12'd1294: rd_data_0 <= 24'h7f0080;
		12'd1295: rd_data_0 <= 24'h7f0080;
		12'd1296: rd_data_0 <= 24'h79007b;
		12'd1297: rd_data_0 <= 24'h810684;
		12'd1298: rd_data_0 <= 24'h78017e;
		12'd1299: rd_data_0 <= 24'h7b0180;
		12'd1300: rd_data_0 <= 24'h79007d;
		12'd1301: rd_data_0 <= 24'h7e0281;
		12'd1302: rd_data_0 <= 24'h77017c;
		12'd1303: rd_data_0 <= 24'h7a017e;
		12'd1304: rd_data_0 <= 24'h830484;
		12'd1305: rd_data_0 <= 24'h860583;
		12'd1306: rd_data_0 <= 24'h840580;
		12'd1307: rd_data_0 <= 24'h780676;
		12'd1308: rd_data_0 <= 24'h630e64;
		12'd1309: rd_data_0 <= 24'h653267;
		12'd1310: rd_data_0 <= 24'h625061;
		12'd1311: rd_data_0 <= 24'h7c8779;
		12'd1312: rd_data_0 <= 24'h9db9a2;
		12'd1313: rd_data_0 <= 24'h97baa3;
		12'd1314: rd_data_0 <= 24'h93b79c;
		12'd1315: rd_data_0 <= 24'h8bae90;
		12'd1316: rd_data_0 <= 24'h8aaf8a;
		12'd1317: rd_data_0 <= 24'h83aa7e;
		12'd1318: rd_data_0 <= 24'h6f9566;
		12'd1319: rd_data_0 <= 24'h7fa774;
		12'd1320: rd_data_0 <= 24'h77aa6d;
		12'd1321: rd_data_0 <= 24'h558f4d;
		12'd1322: rd_data_0 <= 24'h609461;
		12'd1323: rd_data_0 <= 24'h48644d;
		12'd1324: rd_data_0 <= 24'h635667;
		12'd1325: rd_data_0 <= 24'h40013e;
		12'd1326: rd_data_0 <= 24'h751176;
		12'd1327: rd_data_0 <= 24'h75007c;
		12'd1328: rd_data_0 <= 24'h82068a;
		12'd1329: rd_data_0 <= 24'h7f0180;
		12'd1330: rd_data_0 <= 24'h800180;
		12'd1331: rd_data_0 <= 24'h800180;
		12'd1332: rd_data_0 <= 24'h800180;
		12'd1333: rd_data_0 <= 24'h800180;
		12'd1334: rd_data_0 <= 24'h800180;
		12'd1335: rd_data_0 <= 24'h800180;
		12'd1336: rd_data_0 <= 24'h800180;
		12'd1337: rd_data_0 <= 24'h800180;
		12'd1338: rd_data_0 <= 24'h800180;
		12'd1339: rd_data_0 <= 24'h800180;
		12'd1340: rd_data_0 <= 24'h800180;
		12'd1341: rd_data_0 <= 24'h800180;
		12'd1342: rd_data_0 <= 24'h800180;
		12'd1343: rd_data_0 <= 24'h800180;
		12'd1344: rd_data_0 <= 24'h7f007f;
		12'd1345: rd_data_0 <= 24'h7f007f;
		12'd1346: rd_data_0 <= 24'h7f007f;
		12'd1347: rd_data_0 <= 24'h7f007f;
		12'd1348: rd_data_0 <= 24'h7f007f;
		12'd1349: rd_data_0 <= 24'h7f007f;
		12'd1350: rd_data_0 <= 24'h7f007f;
		12'd1351: rd_data_0 <= 24'h7f007f;
		12'd1352: rd_data_0 <= 24'h7f007f;
		12'd1353: rd_data_0 <= 24'h7f007f;
		12'd1354: rd_data_0 <= 24'h7f007f;
		12'd1355: rd_data_0 <= 24'h7f007f;
		12'd1356: rd_data_0 <= 24'h7f007f;
		12'd1357: rd_data_0 <= 24'h7f007f;
		12'd1358: rd_data_0 <= 24'h80007f;
		12'd1359: rd_data_0 <= 24'h7b017e;
		12'd1360: rd_data_0 <= 24'h790d81;
		12'd1361: rd_data_0 <= 24'h721283;
		12'd1362: rd_data_0 <= 24'h620975;
		12'd1363: rd_data_0 <= 24'h6c0d7b;
		12'd1364: rd_data_0 <= 24'h720678;
		12'd1365: rd_data_0 <= 24'h7a057b;
		12'd1366: rd_data_0 <= 24'h790679;
		12'd1367: rd_data_0 <= 24'h7c097d;
		12'd1368: rd_data_0 <= 24'h800b81;
		12'd1369: rd_data_0 <= 24'h810d7e;
		12'd1370: rd_data_0 <= 24'h7c0d74;
		12'd1371: rd_data_0 <= 24'h63095b;
		12'd1372: rd_data_0 <= 24'h5c2f5d;
		12'd1373: rd_data_0 <= 24'h888b90;
		12'd1374: rd_data_0 <= 24'h9dc0a1;
		12'd1375: rd_data_0 <= 24'h99d099;
		12'd1376: rd_data_0 <= 24'h9edea3;
		12'd1377: rd_data_0 <= 24'ha0e1aa;
		12'd1378: rd_data_0 <= 24'ha2e5ac;
		12'd1379: rd_data_0 <= 24'ha2e6a8;
		12'd1380: rd_data_0 <= 24'ha0e4a0;
		12'd1381: rd_data_0 <= 24'ha3e79f;
		12'd1382: rd_data_0 <= 24'h81c679;
		12'd1383: rd_data_0 <= 24'h4c9040;
		12'd1384: rd_data_0 <= 24'h61a458;
		12'd1385: rd_data_0 <= 24'h7cbc7a;
		12'd1386: rd_data_0 <= 24'h72aa75;
		12'd1387: rd_data_0 <= 24'h4b6f52;
		12'd1388: rd_data_0 <= 24'h444248;
		12'd1389: rd_data_0 <= 24'h2e0030;
		12'd1390: rd_data_0 <= 24'h6b0f70;
		12'd1391: rd_data_0 <= 24'h770282;
		12'd1392: rd_data_0 <= 24'h80028b;
		12'd1393: rd_data_0 <= 24'h800083;
		12'd1394: rd_data_0 <= 24'h810180;
		12'd1395: rd_data_0 <= 24'h810180;
		12'd1396: rd_data_0 <= 24'h810180;
		12'd1397: rd_data_0 <= 24'h810180;
		12'd1398: rd_data_0 <= 24'h810180;
		12'd1399: rd_data_0 <= 24'h810180;
		12'd1400: rd_data_0 <= 24'h810180;
		12'd1401: rd_data_0 <= 24'h810180;
		12'd1402: rd_data_0 <= 24'h810180;
		12'd1403: rd_data_0 <= 24'h810180;
		12'd1404: rd_data_0 <= 24'h810180;
		12'd1405: rd_data_0 <= 24'h810180;
		12'd1406: rd_data_0 <= 24'h810180;
		12'd1407: rd_data_0 <= 24'h810180;
		12'd1408: rd_data_0 <= 24'h7f007f;
		12'd1409: rd_data_0 <= 24'h7f007f;
		12'd1410: rd_data_0 <= 24'h7f007f;
		12'd1411: rd_data_0 <= 24'h7f007f;
		12'd1412: rd_data_0 <= 24'h7f007f;
		12'd1413: rd_data_0 <= 24'h7f007f;
		12'd1414: rd_data_0 <= 24'h7f007f;
		12'd1415: rd_data_0 <= 24'h7f007f;
		12'd1416: rd_data_0 <= 24'h7f007f;
		12'd1417: rd_data_0 <= 24'h7f007f;
		12'd1418: rd_data_0 <= 24'h7f007e;
		12'd1419: rd_data_0 <= 24'h7f007e;
		12'd1420: rd_data_0 <= 24'h7e017e;
		12'd1421: rd_data_0 <= 24'h7e017e;
		12'd1422: rd_data_0 <= 24'h80007e;
		12'd1423: rd_data_0 <= 24'h76067c;
		12'd1424: rd_data_0 <= 24'h571171;
		12'd1425: rd_data_0 <= 24'h401667;
		12'd1426: rd_data_0 <= 24'h3d1c69;
		12'd1427: rd_data_0 <= 24'h4a1f70;
		12'd1428: rd_data_0 <= 24'h5f1974;
		12'd1429: rd_data_0 <= 24'h691071;
		12'd1430: rd_data_0 <= 24'h6b0f70;
		12'd1431: rd_data_0 <= 24'h670b6d;
		12'd1432: rd_data_0 <= 24'h650a6a;
		12'd1433: rd_data_0 <= 24'h5d0961;
		12'd1434: rd_data_0 <= 24'h57185d;
		12'd1435: rd_data_0 <= 24'h603c68;
		12'd1436: rd_data_0 <= 24'h8b8b9a;
		12'd1437: rd_data_0 <= 24'habcbbf;
		12'd1438: rd_data_0 <= 24'ha6ddbd;
		12'd1439: rd_data_0 <= 24'h9ee5b8;
		12'd1440: rd_data_0 <= 24'ha4eebd;
		12'd1441: rd_data_0 <= 24'h6ab283;
		12'd1442: rd_data_0 <= 24'h225e2b;
		12'd1443: rd_data_0 <= 24'h3b7a42;
		12'd1444: rd_data_0 <= 24'h5da96c;
		12'd1445: rd_data_0 <= 24'h57a25f;
		12'd1446: rd_data_0 <= 24'h68b36c;
		12'd1447: rd_data_0 <= 24'h73be76;
		12'd1448: rd_data_0 <= 24'h64b46b;
		12'd1449: rd_data_0 <= 24'h71c17e;
		12'd1450: rd_data_0 <= 24'h68ac73;
		12'd1451: rd_data_0 <= 24'h4b7852;
		12'd1452: rd_data_0 <= 24'h303c35;
		12'd1453: rd_data_0 <= 24'h1f0024;
		12'd1454: rd_data_0 <= 24'h681b6c;
		12'd1455: rd_data_0 <= 24'h7e0782;
		12'd1456: rd_data_0 <= 24'h880389;
		12'd1457: rd_data_0 <= 24'h810080;
		12'd1458: rd_data_0 <= 24'h810180;
		12'd1459: rd_data_0 <= 24'h820081;
		12'd1460: rd_data_0 <= 24'h820081;
		12'd1461: rd_data_0 <= 24'h810180;
		12'd1462: rd_data_0 <= 24'h810180;
		12'd1463: rd_data_0 <= 24'h810180;
		12'd1464: rd_data_0 <= 24'h810180;
		12'd1465: rd_data_0 <= 24'h810180;
		12'd1466: rd_data_0 <= 24'h810180;
		12'd1467: rd_data_0 <= 24'h810180;
		12'd1468: rd_data_0 <= 24'h810180;
		12'd1469: rd_data_0 <= 24'h810180;
		12'd1470: rd_data_0 <= 24'h810180;
		12'd1471: rd_data_0 <= 24'h810180;
		12'd1472: rd_data_0 <= 24'h7f007f;
		12'd1473: rd_data_0 <= 24'h7f007f;
		12'd1474: rd_data_0 <= 24'h7f007f;
		12'd1475: rd_data_0 <= 24'h7f007f;
		12'd1476: rd_data_0 <= 24'h7f007f;
		12'd1477: rd_data_0 <= 24'h7f007f;
		12'd1478: rd_data_0 <= 24'h7f007f;
		12'd1479: rd_data_0 <= 24'h7f007f;
		12'd1480: rd_data_0 <= 24'h7f007f;
		12'd1481: rd_data_0 <= 24'h7f007f;
		12'd1482: rd_data_0 <= 24'h7f007d;
		12'd1483: rd_data_0 <= 24'h7f007d;
		12'd1484: rd_data_0 <= 24'h7e017d;
		12'd1485: rd_data_0 <= 24'h7e017d;
		12'd1486: rd_data_0 <= 24'h80007e;
		12'd1487: rd_data_0 <= 24'h6d0576;
		12'd1488: rd_data_0 <= 24'h64408b;
		12'd1489: rd_data_0 <= 24'h808bbb;
		12'd1490: rd_data_0 <= 24'h90a6d0;
		12'd1491: rd_data_0 <= 24'h444f7d;
		12'd1492: rd_data_0 <= 24'h3c2861;
		12'd1493: rd_data_0 <= 24'h4f2363;
		12'd1494: rd_data_0 <= 24'h5f2f71;
		12'd1495: rd_data_0 <= 24'h633577;
		12'd1496: rd_data_0 <= 24'h5e3271;
		12'd1497: rd_data_0 <= 24'h56336b;
		12'd1498: rd_data_0 <= 24'h484163;
		12'd1499: rd_data_0 <= 24'h485d67;
		12'd1500: rd_data_0 <= 24'h5b867d;
		12'd1501: rd_data_0 <= 24'h548f7a;
		12'd1502: rd_data_0 <= 24'h4a9177;
		12'd1503: rd_data_0 <= 24'h38856a;
		12'd1504: rd_data_0 <= 24'h287353;
		12'd1505: rd_data_0 <= 24'h4a9472;
		12'd1506: rd_data_0 <= 24'h67a884;
		12'd1507: rd_data_0 <= 24'h326941;
		12'd1508: rd_data_0 <= 24'h316e3f;
		12'd1509: rd_data_0 <= 24'h74bd86;
		12'd1510: rd_data_0 <= 24'h7ec88c;
		12'd1511: rd_data_0 <= 24'h92df9e;
		12'd1512: rd_data_0 <= 24'h79d18a;
		12'd1513: rd_data_0 <= 24'h62c07b;
		12'd1514: rd_data_0 <= 24'h66b778;
		12'd1515: rd_data_0 <= 24'h599363;
		12'd1516: rd_data_0 <= 24'h3b5a43;
		12'd1517: rd_data_0 <= 24'h45434f;
		12'd1518: rd_data_0 <= 24'h3a073f;
		12'd1519: rd_data_0 <= 24'h760e73;
		12'd1520: rd_data_0 <= 24'h7f007a;
		12'd1521: rd_data_0 <= 24'h820180;
		12'd1522: rd_data_0 <= 24'h810081;
		12'd1523: rd_data_0 <= 24'h820082;
		12'd1524: rd_data_0 <= 24'h820082;
		12'd1525: rd_data_0 <= 24'h810180;
		12'd1526: rd_data_0 <= 24'h810180;
		12'd1527: rd_data_0 <= 24'h810180;
		12'd1528: rd_data_0 <= 24'h810180;
		12'd1529: rd_data_0 <= 24'h810180;
		12'd1530: rd_data_0 <= 24'h810180;
		12'd1531: rd_data_0 <= 24'h810180;
		12'd1532: rd_data_0 <= 24'h810180;
		12'd1533: rd_data_0 <= 24'h810180;
		12'd1534: rd_data_0 <= 24'h810180;
		12'd1535: rd_data_0 <= 24'h810180;
		12'd1536: rd_data_0 <= 24'h7f007f;
		12'd1537: rd_data_0 <= 24'h7f007f;
		12'd1538: rd_data_0 <= 24'h7f007f;
		12'd1539: rd_data_0 <= 24'h7f007f;
		12'd1540: rd_data_0 <= 24'h7f007f;
		12'd1541: rd_data_0 <= 24'h7f007f;
		12'd1542: rd_data_0 <= 24'h7f007e;
		12'd1543: rd_data_0 <= 24'h7f007e;
		12'd1544: rd_data_0 <= 24'h7e017e;
		12'd1545: rd_data_0 <= 24'h7e017e;
		12'd1546: rd_data_0 <= 24'h7f007d;
		12'd1547: rd_data_0 <= 24'h7f007d;
		12'd1548: rd_data_0 <= 24'h7e017d;
		12'd1549: rd_data_0 <= 24'h7f007d;
		12'd1550: rd_data_0 <= 24'h82007e;
		12'd1551: rd_data_0 <= 24'h690571;
		12'd1552: rd_data_0 <= 24'h6a5b92;
		12'd1553: rd_data_0 <= 24'ha1d0e1;
		12'd1554: rd_data_0 <= 24'ha9ecef;
		12'd1555: rd_data_0 <= 24'h84c5c5;
		12'd1556: rd_data_0 <= 24'h436e75;
		12'd1557: rd_data_0 <= 24'h2c4453;
		12'd1558: rd_data_0 <= 24'h73889d;
		12'd1559: rd_data_0 <= 24'h95aec3;
		12'd1560: rd_data_0 <= 24'h91aec1;
		12'd1561: rd_data_0 <= 24'h8db2bf;
		12'd1562: rd_data_0 <= 24'h87bebd;
		12'd1563: rd_data_0 <= 24'h6cb7a7;
		12'd1564: rd_data_0 <= 24'h57ad95;
		12'd1565: rd_data_0 <= 24'h57b397;
		12'd1566: rd_data_0 <= 24'h1f775c;
		12'd1567: rd_data_0 <= 24'h287d63;
		12'd1568: rd_data_0 <= 24'h5fb496;
		12'd1569: rd_data_0 <= 24'h80d1af;
		12'd1570: rd_data_0 <= 24'haeefd3;
		12'd1571: rd_data_0 <= 24'h4f7962;
		12'd1572: rd_data_0 <= 24'h325e3d;
		12'd1573: rd_data_0 <= 24'ha2e3b3;
		12'd1574: rd_data_0 <= 24'h90da9c;
		12'd1575: rd_data_0 <= 24'h8bdd93;
		12'd1576: rd_data_0 <= 24'h7cd68b;
		12'd1577: rd_data_0 <= 24'h63c17a;
		12'd1578: rd_data_0 <= 24'h68c17d;
		12'd1579: rd_data_0 <= 24'h5da86a;
		12'd1580: rd_data_0 <= 24'h347042;
		12'd1581: rd_data_0 <= 24'h59806d;
		12'd1582: rd_data_0 <= 24'h413d4f;
		12'd1583: rd_data_0 <= 24'h420444;
		12'd1584: rd_data_0 <= 24'h750f73;
		12'd1585: rd_data_0 <= 24'h80017f;
		12'd1586: rd_data_0 <= 24'h850085;
		12'd1587: rd_data_0 <= 24'h830083;
		12'd1588: rd_data_0 <= 24'h820082;
		12'd1589: rd_data_0 <= 24'h820081;
		12'd1590: rd_data_0 <= 24'h820081;
		12'd1591: rd_data_0 <= 24'h820081;
		12'd1592: rd_data_0 <= 24'h820081;
		12'd1593: rd_data_0 <= 24'h820081;
		12'd1594: rd_data_0 <= 24'h820081;
		12'd1595: rd_data_0 <= 24'h810180;
		12'd1596: rd_data_0 <= 24'h810180;
		12'd1597: rd_data_0 <= 24'h810180;
		12'd1598: rd_data_0 <= 24'h810180;
		12'd1599: rd_data_0 <= 24'h810180;
		12'd1600: rd_data_0 <= 24'h7f007f;
		12'd1601: rd_data_0 <= 24'h7f007f;
		12'd1602: rd_data_0 <= 24'h7f007f;
		12'd1603: rd_data_0 <= 24'h7f007f;
		12'd1604: rd_data_0 <= 24'h7f007f;
		12'd1605: rd_data_0 <= 24'h7f007f;
		12'd1606: rd_data_0 <= 24'h7f007d;
		12'd1607: rd_data_0 <= 24'h7f007d;
		12'd1608: rd_data_0 <= 24'h7e017d;
		12'd1609: rd_data_0 <= 24'h7e017d;
		12'd1610: rd_data_0 <= 24'h7f007d;
		12'd1611: rd_data_0 <= 24'h7f007d;
		12'd1612: rd_data_0 <= 24'h7f007d;
		12'd1613: rd_data_0 <= 24'h7f007d;
		12'd1614: rd_data_0 <= 24'h83007e;
		12'd1615: rd_data_0 <= 24'h680770;
		12'd1616: rd_data_0 <= 24'h63608a;
		12'd1617: rd_data_0 <= 24'h94dad5;
		12'd1618: rd_data_0 <= 24'h60c0a6;
		12'd1619: rd_data_0 <= 24'h7ae0bd;
		12'd1620: rd_data_0 <= 24'h76ceb0;
		12'd1621: rd_data_0 <= 24'h6bb9a0;
		12'd1622: rd_data_0 <= 24'h87d5c6;
		12'd1623: rd_data_0 <= 24'h9bede2;
		12'd1624: rd_data_0 <= 24'h72c7b9;
		12'd1625: rd_data_0 <= 24'h5cb4a0;
		12'd1626: rd_data_0 <= 24'h59b9a0;
		12'd1627: rd_data_0 <= 24'h71dbbe;
		12'd1628: rd_data_0 <= 24'h71e3c3;
		12'd1629: rd_data_0 <= 24'h63d9b7;
		12'd1630: rd_data_0 <= 24'h50bb9d;
		12'd1631: rd_data_0 <= 24'h6ccbaf;
		12'd1632: rd_data_0 <= 24'h96f7d6;
		12'd1633: rd_data_0 <= 24'h8ae6c2;
		12'd1634: rd_data_0 <= 24'h94d6bd;
		12'd1635: rd_data_0 <= 24'h4a6e5e;
		12'd1636: rd_data_0 <= 24'h3c6048;
		12'd1637: rd_data_0 <= 24'hb1ebc1;
		12'd1638: rd_data_0 <= 24'h8fd798;
		12'd1639: rd_data_0 <= 24'h90e593;
		12'd1640: rd_data_0 <= 24'h80d987;
		12'd1641: rd_data_0 <= 24'h68c078;
		12'd1642: rd_data_0 <= 24'h6dc47e;
		12'd1643: rd_data_0 <= 24'h5aae67;
		12'd1644: rd_data_0 <= 24'h257537;
		12'd1645: rd_data_0 <= 24'h377d51;
		12'd1646: rd_data_0 <= 24'h4f7264;
		12'd1647: rd_data_0 <= 24'h1a0724;
		12'd1648: rd_data_0 <= 24'h651c67;
		12'd1649: rd_data_0 <= 24'h7b037c;
		12'd1650: rd_data_0 <= 24'h860086;
		12'd1651: rd_data_0 <= 24'h830083;
		12'd1652: rd_data_0 <= 24'h820082;
		12'd1653: rd_data_0 <= 24'h820082;
		12'd1654: rd_data_0 <= 24'h820082;
		12'd1655: rd_data_0 <= 24'h820082;
		12'd1656: rd_data_0 <= 24'h820082;
		12'd1657: rd_data_0 <= 24'h820082;
		12'd1658: rd_data_0 <= 24'h820082;
		12'd1659: rd_data_0 <= 24'h810180;
		12'd1660: rd_data_0 <= 24'h810180;
		12'd1661: rd_data_0 <= 24'h810180;
		12'd1662: rd_data_0 <= 24'h810180;
		12'd1663: rd_data_0 <= 24'h810180;
		12'd1664: rd_data_0 <= 24'h7f007f;
		12'd1665: rd_data_0 <= 24'h7f007f;
		12'd1666: rd_data_0 <= 24'h7f007f;
		12'd1667: rd_data_0 <= 24'h7f007f;
		12'd1668: rd_data_0 <= 24'h7f007f;
		12'd1669: rd_data_0 <= 24'h7f007f;
		12'd1670: rd_data_0 <= 24'h7f007d;
		12'd1671: rd_data_0 <= 24'h7f007d;
		12'd1672: rd_data_0 <= 24'h7e017d;
		12'd1673: rd_data_0 <= 24'h7e017d;
		12'd1674: rd_data_0 <= 24'h7f017c;
		12'd1675: rd_data_0 <= 24'h7f007c;
		12'd1676: rd_data_0 <= 24'h7f007c;
		12'd1677: rd_data_0 <= 24'h7f007c;
		12'd1678: rd_data_0 <= 24'h81007d;
		12'd1679: rd_data_0 <= 24'h64096e;
		12'd1680: rd_data_0 <= 24'h666d92;
		12'd1681: rd_data_0 <= 24'h47968b;
		12'd1682: rd_data_0 <= 24'h56bd9c;
		12'd1683: rd_data_0 <= 24'h7ce7be;
		12'd1684: rd_data_0 <= 24'h8ef1ca;
		12'd1685: rd_data_0 <= 24'h90efcc;
		12'd1686: rd_data_0 <= 24'h8cf1d6;
		12'd1687: rd_data_0 <= 24'h65d0b9;
		12'd1688: rd_data_0 <= 24'h40a38c;
		12'd1689: rd_data_0 <= 24'h37937b;
		12'd1690: rd_data_0 <= 24'h2e8c73;
		12'd1691: rd_data_0 <= 24'h63caad;
		12'd1692: rd_data_0 <= 24'h7af2d0;
		12'd1693: rd_data_0 <= 24'h5bdeb9;
		12'd1694: rd_data_0 <= 24'h65ddbc;
		12'd1695: rd_data_0 <= 24'h73dec0;
		12'd1696: rd_data_0 <= 24'h72debc;
		12'd1697: rd_data_0 <= 24'h6fd9b5;
		12'd1698: rd_data_0 <= 24'h74cbb0;
		12'd1699: rd_data_0 <= 24'h5a9a85;
		12'd1700: rd_data_0 <= 24'h2d5c44;
		12'd1701: rd_data_0 <= 24'h64926e;
		12'd1702: rd_data_0 <= 24'h9bdda3;
		12'd1703: rd_data_0 <= 24'h94e898;
		12'd1704: rd_data_0 <= 24'h86db8a;
		12'd1705: rd_data_0 <= 24'h73c17a;
		12'd1706: rd_data_0 <= 24'h75c37f;
		12'd1707: rd_data_0 <= 24'h5db069;
		12'd1708: rd_data_0 <= 24'h2a7e3d;
		12'd1709: rd_data_0 <= 24'h20713d;
		12'd1710: rd_data_0 <= 24'h538a6e;
		12'd1711: rd_data_0 <= 24'h354045;
		12'd1712: rd_data_0 <= 24'h390c40;
		12'd1713: rd_data_0 <= 24'h740a75;
		12'd1714: rd_data_0 <= 24'h820181;
		12'd1715: rd_data_0 <= 24'h820182;
		12'd1716: rd_data_0 <= 24'h820082;
		12'd1717: rd_data_0 <= 24'h820082;
		12'd1718: rd_data_0 <= 24'h820082;
		12'd1719: rd_data_0 <= 24'h820082;
		12'd1720: rd_data_0 <= 24'h820181;
		12'd1721: rd_data_0 <= 24'h810181;
		12'd1722: rd_data_0 <= 24'h810181;
		12'd1723: rd_data_0 <= 24'h810180;
		12'd1724: rd_data_0 <= 24'h810180;
		12'd1725: rd_data_0 <= 24'h810180;
		12'd1726: rd_data_0 <= 24'h810180;
		12'd1727: rd_data_0 <= 24'h810180;
		12'd1728: rd_data_0 <= 24'h7f007f;
		12'd1729: rd_data_0 <= 24'h7f007f;
		12'd1730: rd_data_0 <= 24'h7f007f;
		12'd1731: rd_data_0 <= 24'h7f007f;
		12'd1732: rd_data_0 <= 24'h7f007f;
		12'd1733: rd_data_0 <= 24'h7f007f;
		12'd1734: rd_data_0 <= 24'h7f007d;
		12'd1735: rd_data_0 <= 24'h7f007d;
		12'd1736: rd_data_0 <= 24'h7e017d;
		12'd1737: rd_data_0 <= 24'h7e017d;
		12'd1738: rd_data_0 <= 24'h7d027b;
		12'd1739: rd_data_0 <= 24'h7f017b;
		12'd1740: rd_data_0 <= 24'h80007b;
		12'd1741: rd_data_0 <= 24'h7f017b;
		12'd1742: rd_data_0 <= 24'h7d027c;
		12'd1743: rd_data_0 <= 24'h5e0d6e;
		12'd1744: rd_data_0 <= 24'h536185;
		12'd1745: rd_data_0 <= 24'h4fa397;
		12'd1746: rd_data_0 <= 24'h77dfbf;
		12'd1747: rd_data_0 <= 24'h81e9c2;
		12'd1748: rd_data_0 <= 24'h88e9c4;
		12'd1749: rd_data_0 <= 24'h8fedcb;
		12'd1750: rd_data_0 <= 24'h69d2b6;
		12'd1751: rd_data_0 <= 24'h33a38b;
		12'd1752: rd_data_0 <= 24'h369983;
		12'd1753: rd_data_0 <= 24'h348d76;
		12'd1754: rd_data_0 <= 24'h51a891;
		12'd1755: rd_data_0 <= 24'h7edec5;
		12'd1756: rd_data_0 <= 24'h81f7d6;
		12'd1757: rd_data_0 <= 24'h66ebc5;
		12'd1758: rd_data_0 <= 24'h5dd6b4;
		12'd1759: rd_data_0 <= 24'h67d1b4;
		12'd1760: rd_data_0 <= 24'h6ad8b7;
		12'd1761: rd_data_0 <= 24'h65d8b4;
		12'd1762: rd_data_0 <= 24'h66d3b5;
		12'd1763: rd_data_0 <= 24'h5cbba2;
		12'd1764: rd_data_0 <= 24'h18543b;
		12'd1765: rd_data_0 <= 24'h345738;
		12'd1766: rd_data_0 <= 24'ha7e5b0;
		12'd1767: rd_data_0 <= 24'h8cde94;
		12'd1768: rd_data_0 <= 24'h7ece82;
		12'd1769: rd_data_0 <= 24'h7bc17b;
		12'd1770: rd_data_0 <= 24'h7dc581;
		12'd1771: rd_data_0 <= 24'h63b36e;
		12'd1772: rd_data_0 <= 24'h378949;
		12'd1773: rd_data_0 <= 24'h2b7d45;
		12'd1774: rd_data_0 <= 24'h397b54;
		12'd1775: rd_data_0 <= 24'h456857;
		12'd1776: rd_data_0 <= 24'h14001d;
		12'd1777: rd_data_0 <= 24'h6d156d;
		12'd1778: rd_data_0 <= 24'h7c047a;
		12'd1779: rd_data_0 <= 24'h7f017e;
		12'd1780: rd_data_0 <= 24'h820182;
		12'd1781: rd_data_0 <= 24'h830083;
		12'd1782: rd_data_0 <= 24'h830083;
		12'd1783: rd_data_0 <= 24'h800080;
		12'd1784: rd_data_0 <= 24'h80007f;
		12'd1785: rd_data_0 <= 24'h810180;
		12'd1786: rd_data_0 <= 24'h810180;
		12'd1787: rd_data_0 <= 24'h810180;
		12'd1788: rd_data_0 <= 24'h810180;
		12'd1789: rd_data_0 <= 24'h810180;
		12'd1790: rd_data_0 <= 24'h810180;
		12'd1791: rd_data_0 <= 24'h810180;
		12'd1792: rd_data_0 <= 24'h7f007f;
		12'd1793: rd_data_0 <= 24'h7f007f;
		12'd1794: rd_data_0 <= 24'h7f007f;
		12'd1795: rd_data_0 <= 24'h7f007f;
		12'd1796: rd_data_0 <= 24'h7f007f;
		12'd1797: rd_data_0 <= 24'h7f007f;
		12'd1798: rd_data_0 <= 24'h7f007d;
		12'd1799: rd_data_0 <= 24'h7f007d;
		12'd1800: rd_data_0 <= 24'h7e017d;
		12'd1801: rd_data_0 <= 24'h7d027d;
		12'd1802: rd_data_0 <= 24'h7b037b;
		12'd1803: rd_data_0 <= 24'h7d027b;
		12'd1804: rd_data_0 <= 24'h80007a;
		12'd1805: rd_data_0 <= 24'h7e007a;
		12'd1806: rd_data_0 <= 24'h79057d;
		12'd1807: rd_data_0 <= 24'h530e6a;
		12'd1808: rd_data_0 <= 24'h3e5273;
		12'd1809: rd_data_0 <= 24'h75cdbf;
		12'd1810: rd_data_0 <= 24'h82f0cd;
		12'd1811: rd_data_0 <= 24'h7febc3;
		12'd1812: rd_data_0 <= 24'h8feec9;
		12'd1813: rd_data_0 <= 24'h93eacb;
		12'd1814: rd_data_0 <= 24'h4eab94;
		12'd1815: rd_data_0 <= 24'h2a8d79;
		12'd1816: rd_data_0 <= 24'h2f927c;
		12'd1817: rd_data_0 <= 24'h4fb198;
		12'd1818: rd_data_0 <= 24'h79dcc1;
		12'd1819: rd_data_0 <= 24'h8bf1d5;
		12'd1820: rd_data_0 <= 24'h84f7d7;
		12'd1821: rd_data_0 <= 24'h76efcd;
		12'd1822: rd_data_0 <= 24'h59c4a6;
		12'd1823: rd_data_0 <= 24'h45a188;
		12'd1824: rd_data_0 <= 24'h5dbfa4;
		12'd1825: rd_data_0 <= 24'h69d7ba;
		12'd1826: rd_data_0 <= 24'h65d9bd;
		12'd1827: rd_data_0 <= 24'h58c6ac;
		12'd1828: rd_data_0 <= 24'h11533c;
		12'd1829: rd_data_0 <= 24'h406045;
		12'd1830: rd_data_0 <= 24'hace6b8;
		12'd1831: rd_data_0 <= 24'h76c580;
		12'd1832: rd_data_0 <= 24'h76c279;
		12'd1833: rd_data_0 <= 24'h80c47d;
		12'd1834: rd_data_0 <= 24'h7ac07b;
		12'd1835: rd_data_0 <= 24'h53a360;
		12'd1836: rd_data_0 <= 24'h3e9151;
		12'd1837: rd_data_0 <= 24'h34844b;
		12'd1838: rd_data_0 <= 24'h226e3a;
		12'd1839: rd_data_0 <= 24'h48835a;
		12'd1840: rd_data_0 <= 24'h3d4346;
		12'd1841: rd_data_0 <= 24'h4b0a4a;
		12'd1842: rd_data_0 <= 24'h760a73;
		12'd1843: rd_data_0 <= 24'h7a0379;
		12'd1844: rd_data_0 <= 24'h7f007f;
		12'd1845: rd_data_0 <= 24'h830083;
		12'd1846: rd_data_0 <= 24'h830083;
		12'd1847: rd_data_0 <= 24'h7f007f;
		12'd1848: rd_data_0 <= 24'h7f017e;
		12'd1849: rd_data_0 <= 24'h800080;
		12'd1850: rd_data_0 <= 24'h80007f;
		12'd1851: rd_data_0 <= 24'h80007f;
		12'd1852: rd_data_0 <= 24'h80007f;
		12'd1853: rd_data_0 <= 24'h810180;
		12'd1854: rd_data_0 <= 24'h810180;
		12'd1855: rd_data_0 <= 24'h80007f;
		12'd1856: rd_data_0 <= 24'h7f007f;
		12'd1857: rd_data_0 <= 24'h7f007f;
		12'd1858: rd_data_0 <= 24'h7f007f;
		12'd1859: rd_data_0 <= 24'h7f007f;
		12'd1860: rd_data_0 <= 24'h7f007f;
		12'd1861: rd_data_0 <= 24'h7f007f;
		12'd1862: rd_data_0 <= 24'h7f007d;
		12'd1863: rd_data_0 <= 24'h7f007d;
		12'd1864: rd_data_0 <= 24'h7e017d;
		12'd1865: rd_data_0 <= 24'h7c027d;
		12'd1866: rd_data_0 <= 24'h7b037b;
		12'd1867: rd_data_0 <= 24'h7c027b;
		12'd1868: rd_data_0 <= 24'h7c0076;
		12'd1869: rd_data_0 <= 24'h7f027b;
		12'd1870: rd_data_0 <= 24'h71057a;
		12'd1871: rd_data_0 <= 24'h652782;
		12'd1872: rd_data_0 <= 24'h344364;
		12'd1873: rd_data_0 <= 24'h7bc6bb;
		12'd1874: rd_data_0 <= 24'h79e0bf;
		12'd1875: rd_data_0 <= 24'h7de9c1;
		12'd1876: rd_data_0 <= 24'h8cebc6;
		12'd1877: rd_data_0 <= 24'h8de3c5;
		12'd1878: rd_data_0 <= 24'h74c8b4;
		12'd1879: rd_data_0 <= 24'h6dc3b4;
		12'd1880: rd_data_0 <= 24'h63c4af;
		12'd1881: rd_data_0 <= 24'h7ae5c9;
		12'd1882: rd_data_0 <= 24'h86f3d5;
		12'd1883: rd_data_0 <= 24'h77e2c4;
		12'd1884: rd_data_0 <= 24'h8bf0d4;
		12'd1885: rd_data_0 <= 24'h6fc7b0;
		12'd1886: rd_data_0 <= 24'h6db2a2;
		12'd1887: rd_data_0 <= 24'h88c0b4;
		12'd1888: rd_data_0 <= 24'h4d9386;
		12'd1889: rd_data_0 <= 24'h4aa794;
		12'd1890: rd_data_0 <= 24'h63d1bb;
		12'd1891: rd_data_0 <= 24'h42b19b;
		12'd1892: rd_data_0 <= 24'h337f6b;
		12'd1893: rd_data_0 <= 24'h355c47;
		12'd1894: rd_data_0 <= 24'h5d926b;
		12'd1895: rd_data_0 <= 24'h77c485;
		12'd1896: rd_data_0 <= 24'h76c37a;
		12'd1897: rd_data_0 <= 24'h72b970;
		12'd1898: rd_data_0 <= 24'h53a057;
		12'd1899: rd_data_0 <= 24'h419653;
		12'd1900: rd_data_0 <= 24'h3c8f51;
		12'd1901: rd_data_0 <= 24'h37854a;
		12'd1902: rd_data_0 <= 24'h257537;
		12'd1903: rd_data_0 <= 24'h4e9a5d;
		12'd1904: rd_data_0 <= 24'h526b59;
		12'd1905: rd_data_0 <= 24'h30002d;
		12'd1906: rd_data_0 <= 24'h700f6b;
		12'd1907: rd_data_0 <= 24'h770575;
		12'd1908: rd_data_0 <= 24'h7c007d;
		12'd1909: rd_data_0 <= 24'h840084;
		12'd1910: rd_data_0 <= 24'h820083;
		12'd1911: rd_data_0 <= 24'h7d007d;
		12'd1912: rd_data_0 <= 24'h7c017b;
		12'd1913: rd_data_0 <= 24'h7e007e;
		12'd1914: rd_data_0 <= 24'h7f007f;
		12'd1915: rd_data_0 <= 24'h7f007f;
		12'd1916: rd_data_0 <= 24'h7f007f;
		12'd1917: rd_data_0 <= 24'h810180;
		12'd1918: rd_data_0 <= 24'h810180;
		12'd1919: rd_data_0 <= 24'h7f007f;
		12'd1920: rd_data_0 <= 24'h7f007f;
		12'd1921: rd_data_0 <= 24'h7f007f;
		12'd1922: rd_data_0 <= 24'h7f007f;
		12'd1923: rd_data_0 <= 24'h7f007f;
		12'd1924: rd_data_0 <= 24'h7f007f;
		12'd1925: rd_data_0 <= 24'h7f007f;
		12'd1926: rd_data_0 <= 24'h7f007d;
		12'd1927: rd_data_0 <= 24'h7f007d;
		12'd1928: rd_data_0 <= 24'h7e017d;
		12'd1929: rd_data_0 <= 24'h7c027d;
		12'd1930: rd_data_0 <= 24'h7a037c;
		12'd1931: rd_data_0 <= 24'h7b037c;
		12'd1932: rd_data_0 <= 24'h7f0079;
		12'd1933: rd_data_0 <= 24'h80037d;
		12'd1934: rd_data_0 <= 24'h6a0579;
		12'd1935: rd_data_0 <= 24'h672883;
		12'd1936: rd_data_0 <= 24'h4e3f69;
		12'd1937: rd_data_0 <= 24'h769697;
		12'd1938: rd_data_0 <= 24'h80cab2;
		12'd1939: rd_data_0 <= 24'h78dab4;
		12'd1940: rd_data_0 <= 24'h86e7c2;
		12'd1941: rd_data_0 <= 24'h8ae6c8;
		12'd1942: rd_data_0 <= 24'h96edd9;
		12'd1943: rd_data_0 <= 24'h7dd1c5;
		12'd1944: rd_data_0 <= 24'h5cbaa6;
		12'd1945: rd_data_0 <= 24'h72dabf;
		12'd1946: rd_data_0 <= 24'h76e3c5;
		12'd1947: rd_data_0 <= 24'h7bdcc3;
		12'd1948: rd_data_0 <= 24'h7db9ac;
		12'd1949: rd_data_0 <= 24'h5f7374;
		12'd1950: rd_data_0 <= 24'h6b656e;
		12'd1951: rd_data_0 <= 24'hc4bdc7;
		12'd1952: rd_data_0 <= 24'hacc6c8;
		12'd1953: rd_data_0 <= 24'h498a86;
		12'd1954: rd_data_0 <= 24'h389287;
		12'd1955: rd_data_0 <= 24'h339386;
		12'd1956: rd_data_0 <= 24'h499588;
		12'd1957: rd_data_0 <= 24'h305a4a;
		12'd1958: rd_data_0 <= 24'h0a3613;
		12'd1959: rd_data_0 <= 24'h539e63;
		12'd1960: rd_data_0 <= 24'h5ead65;
		12'd1961: rd_data_0 <= 24'h4fa151;
		12'd1962: rd_data_0 <= 24'h3c9748;
		12'd1963: rd_data_0 <= 24'h36954f;
		12'd1964: rd_data_0 <= 24'h368d4f;
		12'd1965: rd_data_0 <= 24'h3f8a4e;
		12'd1966: rd_data_0 <= 24'h23702c;
		12'd1967: rd_data_0 <= 24'h47984d;
		12'd1968: rd_data_0 <= 24'h466947;
		12'd1969: rd_data_0 <= 24'h2c0224;
		12'd1970: rd_data_0 <= 24'h6a1365;
		12'd1971: rd_data_0 <= 24'h740573;
		12'd1972: rd_data_0 <= 24'h7b007e;
		12'd1973: rd_data_0 <= 24'h840086;
		12'd1974: rd_data_0 <= 24'h820083;
		12'd1975: rd_data_0 <= 24'h7c007b;
		12'd1976: rd_data_0 <= 24'h7b017a;
		12'd1977: rd_data_0 <= 24'h7e017d;
		12'd1978: rd_data_0 <= 24'h7f007f;
		12'd1979: rd_data_0 <= 24'h7f007f;
		12'd1980: rd_data_0 <= 24'h7f007f;
		12'd1981: rd_data_0 <= 24'h810180;
		12'd1982: rd_data_0 <= 24'h810180;
		12'd1983: rd_data_0 <= 24'h7f007f;
		12'd1984: rd_data_0 <= 24'h7f007f;
		12'd1985: rd_data_0 <= 24'h7f007f;
		12'd1986: rd_data_0 <= 24'h7f007f;
		12'd1987: rd_data_0 <= 24'h7f007f;
		12'd1988: rd_data_0 <= 24'h7f007f;
		12'd1989: rd_data_0 <= 24'h7f007f;
		12'd1990: rd_data_0 <= 24'h7f007d;
		12'd1991: rd_data_0 <= 24'h7f007d;
		12'd1992: rd_data_0 <= 24'h7e017d;
		12'd1993: rd_data_0 <= 24'h7c027d;
		12'd1994: rd_data_0 <= 24'h7a037d;
		12'd1995: rd_data_0 <= 24'h7b037d;
		12'd1996: rd_data_0 <= 24'h80007a;
		12'd1997: rd_data_0 <= 24'h7b0379;
		12'd1998: rd_data_0 <= 24'h630c76;
		12'd1999: rd_data_0 <= 24'h4d1365;
		12'd2000: rd_data_0 <= 24'h6c406e;
		12'd2001: rd_data_0 <= 24'h72616f;
		12'd2002: rd_data_0 <= 24'h9dc8b9;
		12'd2003: rd_data_0 <= 24'h80d8b6;
		12'd2004: rd_data_0 <= 24'h81e6c1;
		12'd2005: rd_data_0 <= 24'h89efcf;
		12'd2006: rd_data_0 <= 24'h71cdba;
		12'd2007: rd_data_0 <= 24'h449a8e;
		12'd2008: rd_data_0 <= 24'h27826f;
		12'd2009: rd_data_0 <= 24'h62c5ab;
		12'd2010: rd_data_0 <= 24'h6fd6b9;
		12'd2011: rd_data_0 <= 24'h91e3cf;
		12'd2012: rd_data_0 <= 24'h829496;
		12'd2013: rd_data_0 <= 24'h703f57;
		12'd2014: rd_data_0 <= 24'h6d1739;
		12'd2015: rd_data_0 <= 24'hbe85a4;
		12'd2016: rd_data_0 <= 24'hffffff;
		12'd2017: rd_data_0 <= 24'h759a9d;
		12'd2018: rd_data_0 <= 24'h135b5b;
		12'd2019: rd_data_0 <= 24'h429490;
		12'd2020: rd_data_0 <= 24'h428b85;
		12'd2021: rd_data_0 <= 24'h2e5c51;
		12'd2022: rd_data_0 <= 24'h00270c;
		12'd2023: rd_data_0 <= 24'h236c3b;
		12'd2024: rd_data_0 <= 24'h479956;
		12'd2025: rd_data_0 <= 24'h399344;
		12'd2026: rd_data_0 <= 24'h399a4c;
		12'd2027: rd_data_0 <= 24'h31924d;
		12'd2028: rd_data_0 <= 24'h378e4e;
		12'd2029: rd_data_0 <= 24'h388043;
		12'd2030: rd_data_0 <= 24'h358138;
		12'd2031: rd_data_0 <= 24'h469544;
		12'd2032: rd_data_0 <= 24'h496c45;
		12'd2033: rd_data_0 <= 24'h2a0322;
		12'd2034: rd_data_0 <= 24'h6a1464;
		12'd2035: rd_data_0 <= 24'h730573;
		12'd2036: rd_data_0 <= 24'h7c007e;
		12'd2037: rd_data_0 <= 24'h840086;
		12'd2038: rd_data_0 <= 24'h820083;
		12'd2039: rd_data_0 <= 24'h7c007b;
		12'd2040: rd_data_0 <= 24'h7b017a;
		12'd2041: rd_data_0 <= 24'h7e017d;
		12'd2042: rd_data_0 <= 24'h7f007f;
		12'd2043: rd_data_0 <= 24'h7f007f;
		12'd2044: rd_data_0 <= 24'h7f007f;
		12'd2045: rd_data_0 <= 24'h810180;
		12'd2046: rd_data_0 <= 24'h810180;
		12'd2047: rd_data_0 <= 24'h7f007f;

        endcase

        case (i_rd_addr)
		12'd0000: rd_data_1 <= 24'h7f007f;
		12'd0001: rd_data_1 <= 24'h7f007f;
		12'd0002: rd_data_1 <= 24'h7f007f;
		12'd0003: rd_data_1 <= 24'h7f007f;
		12'd0004: rd_data_1 <= 24'h7f007f;
		12'd0005: rd_data_1 <= 24'h7f007f;
		12'd0006: rd_data_1 <= 24'h7f007e;
		12'd0007: rd_data_1 <= 24'h7f007e;
		12'd0008: rd_data_1 <= 24'h7d017e;
		12'd0009: rd_data_1 <= 24'h7c027e;
		12'd0010: rd_data_1 <= 24'h7c027e;
		12'd0011: rd_data_1 <= 24'h7d027d;
		12'd0012: rd_data_1 <= 24'h7d0078;
		12'd0013: rd_data_1 <= 24'h700572;
		12'd0014: rd_data_1 <= 24'h612a74;
		12'd0015: rd_data_1 <= 24'h88699a;
		12'd0016: rd_data_1 <= 24'h864e72;
		12'd0017: rd_data_1 <= 24'hbc98ac;
		12'd0018: rd_data_1 <= 24'h98b4ab;
		12'd0019: rd_data_1 <= 24'h7ccfb2;
		12'd0020: rd_data_1 <= 24'h82eac8;
		12'd0021: rd_data_1 <= 24'h8bf6d8;
		12'd0022: rd_data_1 <= 24'h4eab9b;
		12'd0023: rd_data_1 <= 24'h308479;
		12'd0024: rd_data_1 <= 24'h48a48e;
		12'd0025: rd_data_1 <= 24'h79ddbd;
		12'd0026: rd_data_1 <= 24'h83e6c9;
		12'd0027: rd_data_1 <= 24'h86c8bb;
		12'd0028: rd_data_1 <= 24'h847584;
		12'd0029: rd_data_1 <= 24'hb07095;
		12'd0030: rd_data_1 <= 24'haa3c69;
		12'd0031: rd_data_1 <= 24'h9b3657;
		12'd0032: rd_data_1 <= 24'he1c2cc;
		12'd0033: rd_data_1 <= 24'hbbd2d5;
		12'd0034: rd_data_1 <= 24'h468a8f;
		12'd0035: rd_data_1 <= 24'h3d9793;
		12'd0036: rd_data_1 <= 24'h439892;
		12'd0037: rd_data_1 <= 24'h286860;
		12'd0038: rd_data_1 <= 24'h0e4839;
		12'd0039: rd_data_1 <= 24'h276f54;
		12'd0040: rd_data_1 <= 24'h2b7e4d;
		12'd0041: rd_data_1 <= 24'h3c9655;
		12'd0042: rd_data_1 <= 24'h358f4d;
		12'd0043: rd_data_1 <= 24'h3d9254;
		12'd0044: rd_data_1 <= 24'h408f52;
		12'd0045: rd_data_1 <= 24'h236d2e;
		12'd0046: rd_data_1 <= 24'h46924b;
		12'd0047: rd_data_1 <= 24'h4f974f;
		12'd0048: rd_data_1 <= 24'h526750;
		12'd0049: rd_data_1 <= 24'h34002f;
		12'd0050: rd_data_1 <= 24'h720c6f;
		12'd0051: rd_data_1 <= 24'h7c097b;
		12'd0052: rd_data_1 <= 24'h7a007b;
		12'd0053: rd_data_1 <= 24'h820084;
		12'd0054: rd_data_1 <= 24'h810082;
		12'd0055: rd_data_1 <= 24'h7d007c;
		12'd0056: rd_data_1 <= 24'h7b017b;
		12'd0057: rd_data_1 <= 24'h7e017e;
		12'd0058: rd_data_1 <= 24'h7f007f;
		12'd0059: rd_data_1 <= 24'h7f007f;
		12'd0060: rd_data_1 <= 24'h7f007f;
		12'd0061: rd_data_1 <= 24'h800180;
		12'd0062: rd_data_1 <= 24'h800180;
		12'd0063: rd_data_1 <= 24'h7f007f;
		12'd0064: rd_data_1 <= 24'h7f007f;
		12'd0065: rd_data_1 <= 24'h7f007f;
		12'd0066: rd_data_1 <= 24'h7f007f;
		12'd0067: rd_data_1 <= 24'h7f007f;
		12'd0068: rd_data_1 <= 24'h7f007f;
		12'd0069: rd_data_1 <= 24'h7f007f;
		12'd0070: rd_data_1 <= 24'h7f007f;
		12'd0071: rd_data_1 <= 24'h7e007f;
		12'd0072: rd_data_1 <= 24'h7b027f;
		12'd0073: rd_data_1 <= 24'h7b027f;
		12'd0074: rd_data_1 <= 24'h7c017f;
		12'd0075: rd_data_1 <= 24'h7e007f;
		12'd0076: rd_data_1 <= 24'h7d007c;
		12'd0077: rd_data_1 <= 24'h65036a;
		12'd0078: rd_data_1 <= 24'h59436f;
		12'd0079: rd_data_1 <= 24'hdddfeb;
		12'd0080: rd_data_1 <= 24'h89556a;
		12'd0081: rd_data_1 <= 24'hf8d6eb;
		12'd0082: rd_data_1 <= 24'h88a29b;
		12'd0083: rd_data_1 <= 24'h6ec2a6;
		12'd0084: rd_data_1 <= 24'h83f0cf;
		12'd0085: rd_data_1 <= 24'h88f7dc;
		12'd0086: rd_data_1 <= 24'h6ecdbe;
		12'd0087: rd_data_1 <= 24'h61b6ac;
		12'd0088: rd_data_1 <= 24'h7fe1c7;
		12'd0089: rd_data_1 <= 24'h8bf4d1;
		12'd0090: rd_data_1 <= 24'h89e8ce;
		12'd0091: rd_data_1 <= 24'h6fa9a2;
		12'd0092: rd_data_1 <= 24'h604559;
		12'd0093: rd_data_1 <= 24'hd0a3c8;
		12'd0094: rd_data_1 <= 24'hf19ac2;
		12'd0095: rd_data_1 <= 24'ha82744;
		12'd0096: rd_data_1 <= 24'hd495aa;
		12'd0097: rd_data_1 <= 24'hf0ffff;
		12'd0098: rd_data_1 <= 24'h7dc1c6;
		12'd0099: rd_data_1 <= 24'h2d918a;
		12'd0100: rd_data_1 <= 24'h3c9d93;
		12'd0101: rd_data_1 <= 24'h2f807a;
		12'd0102: rd_data_1 <= 24'h2b7470;
		12'd0103: rd_data_1 <= 24'h3f8881;
		12'd0104: rd_data_1 <= 24'h1b6a51;
		12'd0105: rd_data_1 <= 24'h257c50;
		12'd0106: rd_data_1 <= 24'h469766;
		12'd0107: rd_data_1 <= 24'h418958;
		12'd0108: rd_data_1 <= 24'h347c47;
		12'd0109: rd_data_1 <= 24'h2e7a3d;
		12'd0110: rd_data_1 <= 24'h489150;
		12'd0111: rd_data_1 <= 24'h487f4a;
		12'd0112: rd_data_1 <= 24'h393539;
		12'd0113: rd_data_1 <= 24'h540653;
		12'd0114: rd_data_1 <= 24'h7d047c;
		12'd0115: rd_data_1 <= 24'h820a82;
		12'd0116: rd_data_1 <= 24'h7a017b;
		12'd0117: rd_data_1 <= 24'h7e0080;
		12'd0118: rd_data_1 <= 24'h7e0080;
		12'd0119: rd_data_1 <= 24'h7d027d;
		12'd0120: rd_data_1 <= 24'h7c027d;
		12'd0121: rd_data_1 <= 24'h7e007f;
		12'd0122: rd_data_1 <= 24'h7e007f;
		12'd0123: rd_data_1 <= 24'h7e007f;
		12'd0124: rd_data_1 <= 24'h7e007f;
		12'd0125: rd_data_1 <= 24'h7f007f;
		12'd0126: rd_data_1 <= 24'h7f007f;
		12'd0127: rd_data_1 <= 24'h7f007f;
		12'd0128: rd_data_1 <= 24'h7f007f;
		12'd0129: rd_data_1 <= 24'h7f007f;
		12'd0130: rd_data_1 <= 24'h7f007f;
		12'd0131: rd_data_1 <= 24'h7f007f;
		12'd0132: rd_data_1 <= 24'h7f007f;
		12'd0133: rd_data_1 <= 24'h7f007f;
		12'd0134: rd_data_1 <= 24'h7f007f;
		12'd0135: rd_data_1 <= 24'h7e007f;
		12'd0136: rd_data_1 <= 24'h7b0280;
		12'd0137: rd_data_1 <= 24'h7b0280;
		12'd0138: rd_data_1 <= 24'h7c017f;
		12'd0139: rd_data_1 <= 24'h7d017f;
		12'd0140: rd_data_1 <= 24'h7c007c;
		12'd0141: rd_data_1 <= 24'h67086e;
		12'd0142: rd_data_1 <= 24'h534871;
		12'd0143: rd_data_1 <= 24'hcce0e5;
		12'd0144: rd_data_1 <= 24'h674553;
		12'd0145: rd_data_1 <= 24'h90707f;
		12'd0146: rd_data_1 <= 24'h61897d;
		12'd0147: rd_data_1 <= 24'h5cc2a2;
		12'd0148: rd_data_1 <= 24'h6be3c1;
		12'd0149: rd_data_1 <= 24'h6ee3c7;
		12'd0150: rd_data_1 <= 24'h78e2cf;
		12'd0151: rd_data_1 <= 24'h7de3d1;
		12'd0152: rd_data_1 <= 24'h77e5ca;
		12'd0153: rd_data_1 <= 24'h70e2c1;
		12'd0154: rd_data_1 <= 24'h70d8bf;
		12'd0155: rd_data_1 <= 24'h62a89e;
		12'd0156: rd_data_1 <= 24'h43434e;
		12'd0157: rd_data_1 <= 24'h7b576d;
		12'd0158: rd_data_1 <= 24'hce8fa2;
		12'd0159: rd_data_1 <= 24'hd17e8c;
		12'd0160: rd_data_1 <= 24'hd9b7c3;
		12'd0161: rd_data_1 <= 24'hc1d9e2;
		12'd0162: rd_data_1 <= 24'h67a7ac;
		12'd0163: rd_data_1 <= 24'h3c9692;
		12'd0164: rd_data_1 <= 24'h38988f;
		12'd0165: rd_data_1 <= 24'h39948d;
		12'd0166: rd_data_1 <= 24'h3a8989;
		12'd0167: rd_data_1 <= 24'h4c9394;
		12'd0168: rd_data_1 <= 24'h3a857e;
		12'd0169: rd_data_1 <= 24'h1a6c5b;
		12'd0170: rd_data_1 <= 24'h24745c;
		12'd0171: rd_data_1 <= 24'h257053;
		12'd0172: rd_data_1 <= 24'h348254;
		12'd0173: rd_data_1 <= 24'h489858;
		12'd0174: rd_data_1 <= 24'h519055;
		12'd0175: rd_data_1 <= 24'h496248;
		12'd0176: rd_data_1 <= 24'h1f001d;
		12'd0177: rd_data_1 <= 24'h761377;
		12'd0178: rd_data_1 <= 24'h820482;
		12'd0179: rd_data_1 <= 24'h80057f;
		12'd0180: rd_data_1 <= 24'h7f0480;
		12'd0181: rd_data_1 <= 24'h7e007f;
		12'd0182: rd_data_1 <= 24'h7e007f;
		12'd0183: rd_data_1 <= 24'h7d017e;
		12'd0184: rd_data_1 <= 24'h7d017e;
		12'd0185: rd_data_1 <= 24'h7e007f;
		12'd0186: rd_data_1 <= 24'h7e007f;
		12'd0187: rd_data_1 <= 24'h7e007f;
		12'd0188: rd_data_1 <= 24'h7e007f;
		12'd0189: rd_data_1 <= 24'h7f007f;
		12'd0190: rd_data_1 <= 24'h7f007f;
		12'd0191: rd_data_1 <= 24'h7f007f;
		12'd0192: rd_data_1 <= 24'h7f007f;
		12'd0193: rd_data_1 <= 24'h7f007f;
		12'd0194: rd_data_1 <= 24'h7f007f;
		12'd0195: rd_data_1 <= 24'h7f007f;
		12'd0196: rd_data_1 <= 24'h7f007f;
		12'd0197: rd_data_1 <= 24'h7f007f;
		12'd0198: rd_data_1 <= 24'h7f007f;
		12'd0199: rd_data_1 <= 24'h7e0080;
		12'd0200: rd_data_1 <= 24'h7d0082;
		12'd0201: rd_data_1 <= 24'h7b0282;
		12'd0202: rd_data_1 <= 24'h7a037f;
		12'd0203: rd_data_1 <= 24'h7a027f;
		12'd0204: rd_data_1 <= 24'h7f007c;
		12'd0205: rd_data_1 <= 24'h721079;
		12'd0206: rd_data_1 <= 24'h514275;
		12'd0207: rd_data_1 <= 24'h4c6473;
		12'd0208: rd_data_1 <= 24'h786d7a;
		12'd0209: rd_data_1 <= 24'h6c5c62;
		12'd0210: rd_data_1 <= 24'h5e9283;
		12'd0211: rd_data_1 <= 24'h61ccad;
		12'd0212: rd_data_1 <= 24'h60d8b8;
		12'd0213: rd_data_1 <= 24'h5bd4b7;
		12'd0214: rd_data_1 <= 24'h5dd3b9;
		12'd0215: rd_data_1 <= 24'h64d6bf;
		12'd0216: rd_data_1 <= 24'h5bd2b9;
		12'd0217: rd_data_1 <= 24'h5bd1b6;
		12'd0218: rd_data_1 <= 24'h66d4bc;
		12'd0219: rd_data_1 <= 24'h68bdad;
		12'd0220: rd_data_1 <= 24'h618581;
		12'd0221: rd_data_1 <= 24'h675d5f;
		12'd0222: rd_data_1 <= 24'h947d79;
		12'd0223: rd_data_1 <= 24'hada296;
		12'd0224: rd_data_1 <= 24'ha0adaa;
		12'd0225: rd_data_1 <= 24'h79a1a9;
		12'd0226: rd_data_1 <= 24'h417e83;
		12'd0227: rd_data_1 <= 24'h368281;
		12'd0228: rd_data_1 <= 24'h3f9893;
		12'd0229: rd_data_1 <= 24'h399891;
		12'd0230: rd_data_1 <= 24'h409491;
		12'd0231: rd_data_1 <= 24'h4b9092;
		12'd0232: rd_data_1 <= 24'h4e9699;
		12'd0233: rd_data_1 <= 24'h3f8c90;
		12'd0234: rd_data_1 <= 24'h1e6e6d;
		12'd0235: rd_data_1 <= 24'h1e7164;
		12'd0236: rd_data_1 <= 24'h2e835d;
		12'd0237: rd_data_1 <= 24'h51a162;
		12'd0238: rd_data_1 <= 24'h538054;
		12'd0239: rd_data_1 <= 24'h3d313a;
		12'd0240: rd_data_1 <= 24'h4e104a;
		12'd0241: rd_data_1 <= 24'h770d77;
		12'd0242: rd_data_1 <= 24'h800481;
		12'd0243: rd_data_1 <= 24'h800581;
		12'd0244: rd_data_1 <= 24'h7f0481;
		12'd0245: rd_data_1 <= 24'h7e007f;
		12'd0246: rd_data_1 <= 24'h7e007f;
		12'd0247: rd_data_1 <= 24'h7e007f;
		12'd0248: rd_data_1 <= 24'h7e007f;
		12'd0249: rd_data_1 <= 24'h7e007f;
		12'd0250: rd_data_1 <= 24'h7e007f;
		12'd0251: rd_data_1 <= 24'h7e007f;
		12'd0252: rd_data_1 <= 24'h7e007f;
		12'd0253: rd_data_1 <= 24'h7f007f;
		12'd0254: rd_data_1 <= 24'h7f007f;
		12'd0255: rd_data_1 <= 24'h7f007f;
		12'd0256: rd_data_1 <= 24'h7f007f;
		12'd0257: rd_data_1 <= 24'h7f007f;
		12'd0258: rd_data_1 <= 24'h7f007f;
		12'd0259: rd_data_1 <= 24'h7f007f;
		12'd0260: rd_data_1 <= 24'h7f007f;
		12'd0261: rd_data_1 <= 24'h7f007f;
		12'd0262: rd_data_1 <= 24'h7f007f;
		12'd0263: rd_data_1 <= 24'h7f0081;
		12'd0264: rd_data_1 <= 24'h7e0084;
		12'd0265: rd_data_1 <= 24'h7d0184;
		12'd0266: rd_data_1 <= 24'h79037f;
		12'd0267: rd_data_1 <= 24'h7a027e;
		12'd0268: rd_data_1 <= 24'h80017f;
		12'd0269: rd_data_1 <= 24'h720a7a;
		12'd0270: rd_data_1 <= 24'h47276a;
		12'd0271: rd_data_1 <= 24'h263150;
		12'd0272: rd_data_1 <= 24'h596271;
		12'd0273: rd_data_1 <= 24'h6c757b;
		12'd0274: rd_data_1 <= 24'h99b5b4;
		12'd0275: rd_data_1 <= 24'h9dd3c8;
		12'd0276: rd_data_1 <= 24'h65bca7;
		12'd0277: rd_data_1 <= 24'h5cccb0;
		12'd0278: rd_data_1 <= 24'h68dbbf;
		12'd0279: rd_data_1 <= 24'h48b89e;
		12'd0280: rd_data_1 <= 24'h4fc0a6;
		12'd0281: rd_data_1 <= 24'h6ad9bf;
		12'd0282: rd_data_1 <= 24'h72d7bf;
		12'd0283: rd_data_1 <= 24'h80d2be;
		12'd0284: rd_data_1 <= 24'h98cabb;
		12'd0285: rd_data_1 <= 24'hb3cfc3;
		12'd0286: rd_data_1 <= 24'h90ac9a;
		12'd0287: rd_data_1 <= 24'h628773;
		12'd0288: rd_data_1 <= 24'h436a61;
		12'd0289: rd_data_1 <= 24'h2e5054;
		12'd0290: rd_data_1 <= 24'h285e63;
		12'd0291: rd_data_1 <= 24'h2b7777;
		12'd0292: rd_data_1 <= 24'h388c88;
		12'd0293: rd_data_1 <= 24'h358c88;
		12'd0294: rd_data_1 <= 24'h449693;
		12'd0295: rd_data_1 <= 24'h4a9494;
		12'd0296: rd_data_1 <= 24'h408588;
		12'd0297: rd_data_1 <= 24'h307379;
		12'd0298: rd_data_1 <= 24'h44898e;
		12'd0299: rd_data_1 <= 24'h45918d;
		12'd0300: rd_data_1 <= 24'h1d6951;
		12'd0301: rd_data_1 <= 24'h2f6e43;
		12'd0302: rd_data_1 <= 24'h34453a;
		12'd0303: rd_data_1 <= 24'h3a093d;
		12'd0304: rd_data_1 <= 24'h721671;
		12'd0305: rd_data_1 <= 24'h740173;
		12'd0306: rd_data_1 <= 24'h7e027f;
		12'd0307: rd_data_1 <= 24'h800480;
		12'd0308: rd_data_1 <= 24'h7d017d;
		12'd0309: rd_data_1 <= 24'h7e007f;
		12'd0310: rd_data_1 <= 24'h7e007f;
		12'd0311: rd_data_1 <= 24'h7e007f;
		12'd0312: rd_data_1 <= 24'h7e007f;
		12'd0313: rd_data_1 <= 24'h7e007f;
		12'd0314: rd_data_1 <= 24'h7e007f;
		12'd0315: rd_data_1 <= 24'h7e007f;
		12'd0316: rd_data_1 <= 24'h7e007f;
		12'd0317: rd_data_1 <= 24'h7f007f;
		12'd0318: rd_data_1 <= 24'h7f007f;
		12'd0319: rd_data_1 <= 24'h7f007f;
		12'd0320: rd_data_1 <= 24'h7f007f;
		12'd0321: rd_data_1 <= 24'h7f007f;
		12'd0322: rd_data_1 <= 24'h7f007f;
		12'd0323: rd_data_1 <= 24'h7f007f;
		12'd0324: rd_data_1 <= 24'h7f007f;
		12'd0325: rd_data_1 <= 24'h7f007f;
		12'd0326: rd_data_1 <= 24'h7f007f;
		12'd0327: rd_data_1 <= 24'h800081;
		12'd0328: rd_data_1 <= 24'h810085;
		12'd0329: rd_data_1 <= 24'h7f0086;
		12'd0330: rd_data_1 <= 24'h7a0280;
		12'd0331: rd_data_1 <= 24'h7b037d;
		12'd0332: rd_data_1 <= 24'h7e017d;
		12'd0333: rd_data_1 <= 24'h74077b;
		12'd0334: rd_data_1 <= 24'h4e1368;
		12'd0335: rd_data_1 <= 24'h65578b;
		12'd0336: rd_data_1 <= 24'h2b3a52;
		12'd0337: rd_data_1 <= 24'h5f7478;
		12'd0338: rd_data_1 <= 24'h817b88;
		12'd0339: rd_data_1 <= 24'h837e8b;
		12'd0340: rd_data_1 <= 24'h6d9b93;
		12'd0341: rd_data_1 <= 24'h73c8b1;
		12'd0342: rd_data_1 <= 24'h88ddc7;
		12'd0343: rd_data_1 <= 24'h5daa97;
		12'd0344: rd_data_1 <= 24'h68b5a2;
		12'd0345: rd_data_1 <= 24'h72bca8;
		12'd0346: rd_data_1 <= 24'h609e8c;
		12'd0347: rd_data_1 <= 24'h548775;
		12'd0348: rd_data_1 <= 24'h4f7866;
		12'd0349: rd_data_1 <= 24'h5c7a6a;
		12'd0350: rd_data_1 <= 24'h719d8f;
		12'd0351: rd_data_1 <= 24'h417e72;
		12'd0352: rd_data_1 <= 24'h0d453e;
		12'd0353: rd_data_1 <= 24'h1a3d3f;
		12'd0354: rd_data_1 <= 24'h316668;
		12'd0355: rd_data_1 <= 24'h4d9b9a;
		12'd0356: rd_data_1 <= 24'h2d7c7a;
		12'd0357: rd_data_1 <= 24'h247271;
		12'd0358: rd_data_1 <= 24'h459593;
		12'd0359: rd_data_1 <= 24'h449490;
		12'd0360: rd_data_1 <= 24'h307573;
		12'd0361: rd_data_1 <= 24'h0a4443;
		12'd0362: rd_data_1 <= 24'h1d5858;
		12'd0363: rd_data_1 <= 24'h448584;
		12'd0364: rd_data_1 <= 24'h498a7f;
		12'd0365: rd_data_1 <= 24'h1d4b3a;
		12'd0366: rd_data_1 <= 24'h1f1b30;
		12'd0367: rd_data_1 <= 24'h651c71;
		12'd0368: rd_data_1 <= 24'h6d0073;
		12'd0369: rd_data_1 <= 24'h7c037c;
		12'd0370: rd_data_1 <= 24'h7e017d;
		12'd0371: rd_data_1 <= 24'h7e017d;
		12'd0372: rd_data_1 <= 24'h7e017d;
		12'd0373: rd_data_1 <= 24'h7e007f;
		12'd0374: rd_data_1 <= 24'h7e007f;
		12'd0375: rd_data_1 <= 24'h7e007f;
		12'd0376: rd_data_1 <= 24'h7e007f;
		12'd0377: rd_data_1 <= 24'h7e007f;
		12'd0378: rd_data_1 <= 24'h7e007f;
		12'd0379: rd_data_1 <= 24'h7e007f;
		12'd0380: rd_data_1 <= 24'h7e007f;
		12'd0381: rd_data_1 <= 24'h7f007f;
		12'd0382: rd_data_1 <= 24'h7f007f;
		12'd0383: rd_data_1 <= 24'h7f007f;
		12'd0384: rd_data_1 <= 24'h7f007f;
		12'd0385: rd_data_1 <= 24'h7f007f;
		12'd0386: rd_data_1 <= 24'h7f007f;
		12'd0387: rd_data_1 <= 24'h7f007f;
		12'd0388: rd_data_1 <= 24'h7f007f;
		12'd0389: rd_data_1 <= 24'h7f007f;
		12'd0390: rd_data_1 <= 24'h7f007f;
		12'd0391: rd_data_1 <= 24'h810081;
		12'd0392: rd_data_1 <= 24'h840087;
		12'd0393: rd_data_1 <= 24'h820088;
		12'd0394: rd_data_1 <= 24'h7f0080;
		12'd0395: rd_data_1 <= 24'h7c027c;
		12'd0396: rd_data_1 <= 24'h7c017f;
		12'd0397: rd_data_1 <= 24'h7d0983;
		12'd0398: rd_data_1 <= 24'h650770;
		12'd0399: rd_data_1 <= 24'h4e1361;
		12'd0400: rd_data_1 <= 24'h5a4d78;
		12'd0401: rd_data_1 <= 24'hc7d2dd;
		12'd0402: rd_data_1 <= 24'h6f707e;
		12'd0403: rd_data_1 <= 24'h33323f;
		12'd0404: rd_data_1 <= 24'h5c7373;
		12'd0405: rd_data_1 <= 24'h708c87;
		12'd0406: rd_data_1 <= 24'h828184;
		12'd0407: rd_data_1 <= 24'h9d838f;
		12'd0408: rd_data_1 <= 24'h987b85;
		12'd0409: rd_data_1 <= 24'h71545a;
		12'd0410: rd_data_1 <= 24'h523235;
		12'd0411: rd_data_1 <= 24'h361817;
		12'd0412: rd_data_1 <= 24'h1b0e09;
		12'd0413: rd_data_1 <= 24'h0b0906;
		12'd0414: rd_data_1 <= 24'h608182;
		12'd0415: rd_data_1 <= 24'h71b0b4;
		12'd0416: rd_data_1 <= 24'h3b8283;
		12'd0417: rd_data_1 <= 24'h58999c;
		12'd0418: rd_data_1 <= 24'h5c9b9f;
		12'd0419: rd_data_1 <= 24'h46878a;
		12'd0420: rd_data_1 <= 24'h236d6d;
		12'd0421: rd_data_1 <= 24'h277a77;
		12'd0422: rd_data_1 <= 24'h419690;
		12'd0423: rd_data_1 <= 24'h499a93;
		12'd0424: rd_data_1 <= 24'h448b86;
		12'd0425: rd_data_1 <= 24'h23615b;
		12'd0426: rd_data_1 <= 24'h0b4a46;
		12'd0427: rd_data_1 <= 24'h1b5f5c;
		12'd0428: rd_data_1 <= 24'h559791;
		12'd0429: rd_data_1 <= 24'h50817d;
		12'd0430: rd_data_1 <= 24'h474a65;
		12'd0431: rd_data_1 <= 24'h5a1d6a;
		12'd0432: rd_data_1 <= 24'h68066f;
		12'd0433: rd_data_1 <= 24'h79057a;
		12'd0434: rd_data_1 <= 24'h7e017d;
		12'd0435: rd_data_1 <= 24'h7e017d;
		12'd0436: rd_data_1 <= 24'h7e017d;
		12'd0437: rd_data_1 <= 24'h7e007f;
		12'd0438: rd_data_1 <= 24'h7e007f;
		12'd0439: rd_data_1 <= 24'h7e007f;
		12'd0440: rd_data_1 <= 24'h7e007f;
		12'd0441: rd_data_1 <= 24'h7e007f;
		12'd0442: rd_data_1 <= 24'h7e007f;
		12'd0443: rd_data_1 <= 24'h7e007f;
		12'd0444: rd_data_1 <= 24'h7e007f;
		12'd0445: rd_data_1 <= 24'h7f007f;
		12'd0446: rd_data_1 <= 24'h7f007f;
		12'd0447: rd_data_1 <= 24'h7f007f;
		12'd0448: rd_data_1 <= 24'h7f007f;
		12'd0449: rd_data_1 <= 24'h7f007f;
		12'd0450: rd_data_1 <= 24'h7f007f;
		12'd0451: rd_data_1 <= 24'h7f007f;
		12'd0452: rd_data_1 <= 24'h7f007f;
		12'd0453: rd_data_1 <= 24'h7f007f;
		12'd0454: rd_data_1 <= 24'h7f007f;
		12'd0455: rd_data_1 <= 24'h810082;
		12'd0456: rd_data_1 <= 24'h840089;
		12'd0457: rd_data_1 <= 24'h840088;
		12'd0458: rd_data_1 <= 24'h83007f;
		12'd0459: rd_data_1 <= 24'h80007c;
		12'd0460: rd_data_1 <= 24'h75007a;
		12'd0461: rd_data_1 <= 24'h7b0481;
		12'd0462: rd_data_1 <= 24'h81067e;
		12'd0463: rd_data_1 <= 24'h73096f;
		12'd0464: rd_data_1 <= 24'h571c5e;
		12'd0465: rd_data_1 <= 24'h4f3e63;
		12'd0466: rd_data_1 <= 24'h4a596d;
		12'd0467: rd_data_1 <= 24'h5e757e;
		12'd0468: rd_data_1 <= 24'h4e565e;
		12'd0469: rd_data_1 <= 24'h4c3140;
		12'd0470: rd_data_1 <= 24'h60112e;
		12'd0471: rd_data_1 <= 24'h8b143b;
		12'd0472: rd_data_1 <= 24'ha02348;
		12'd0473: rd_data_1 <= 24'ha72e4c;
		12'd0474: rd_data_1 <= 24'ha9334a;
		12'd0475: rd_data_1 <= 24'ha13b4a;
		12'd0476: rd_data_1 <= 24'h7f3d47;
		12'd0477: rd_data_1 <= 24'h5b474f;
		12'd0478: rd_data_1 <= 24'h45626d;
		12'd0479: rd_data_1 <= 24'h40828f;
		12'd0480: rd_data_1 <= 24'h4d97a2;
		12'd0481: rd_data_1 <= 24'h427f86;
		12'd0482: rd_data_1 <= 24'h38646c;
		12'd0483: rd_data_1 <= 24'h2b5e67;
		12'd0484: rd_data_1 <= 24'h2c7374;
		12'd0485: rd_data_1 <= 24'h429c95;
		12'd0486: rd_data_1 <= 24'h3d968e;
		12'd0487: rd_data_1 <= 24'h44948c;
		12'd0488: rd_data_1 <= 24'h4e9990;
		12'd0489: rd_data_1 <= 24'h358076;
		12'd0490: rd_data_1 <= 24'h1d675e;
		12'd0491: rd_data_1 <= 24'h28746d;
		12'd0492: rd_data_1 <= 24'h4b938f;
		12'd0493: rd_data_1 <= 24'h549294;
		12'd0494: rd_data_1 <= 24'h597387;
		12'd0495: rd_data_1 <= 24'h432759;
		12'd0496: rd_data_1 <= 24'h5d1465;
		12'd0497: rd_data_1 <= 24'h750777;
		12'd0498: rd_data_1 <= 24'h7f017e;
		12'd0499: rd_data_1 <= 24'h7e017d;
		12'd0500: rd_data_1 <= 24'h7e017d;
		12'd0501: rd_data_1 <= 24'h7e007f;
		12'd0502: rd_data_1 <= 24'h7e007f;
		12'd0503: rd_data_1 <= 24'h7e007f;
		12'd0504: rd_data_1 <= 24'h7e007f;
		12'd0505: rd_data_1 <= 24'h7e007f;
		12'd0506: rd_data_1 <= 24'h7e007f;
		12'd0507: rd_data_1 <= 24'h7e007f;
		12'd0508: rd_data_1 <= 24'h7e007f;
		12'd0509: rd_data_1 <= 24'h7f007f;
		12'd0510: rd_data_1 <= 24'h7f007f;
		12'd0511: rd_data_1 <= 24'h7f007f;
		12'd0512: rd_data_1 <= 24'h7f007f;
		12'd0513: rd_data_1 <= 24'h7f007f;
		12'd0514: rd_data_1 <= 24'h7f007f;
		12'd0515: rd_data_1 <= 24'h7f007f;
		12'd0516: rd_data_1 <= 24'h7f007f;
		12'd0517: rd_data_1 <= 24'h7f007f;
		12'd0518: rd_data_1 <= 24'h7f007f;
		12'd0519: rd_data_1 <= 24'h800080;
		12'd0520: rd_data_1 <= 24'h830085;
		12'd0521: rd_data_1 <= 24'h830084;
		12'd0522: rd_data_1 <= 24'h82007e;
		12'd0523: rd_data_1 <= 24'h80007d;
		12'd0524: rd_data_1 <= 24'h75007b;
		12'd0525: rd_data_1 <= 24'h77007c;
		12'd0526: rd_data_1 <= 24'h83007e;
		12'd0527: rd_data_1 <= 24'h7e0075;
		12'd0528: rd_data_1 <= 24'h781675;
		12'd0529: rd_data_1 <= 24'h43054c;
		12'd0530: rd_data_1 <= 24'h1b053a;
		12'd0531: rd_data_1 <= 24'h414267;
		12'd0532: rd_data_1 <= 24'h4f5166;
		12'd0533: rd_data_1 <= 24'h6e6370;
		12'd0534: rd_data_1 <= 24'h724559;
		12'd0535: rd_data_1 <= 24'h914962;
		12'd0536: rd_data_1 <= 24'hc3708c;
		12'd0537: rd_data_1 <= 24'hd27d96;
		12'd0538: rd_data_1 <= 24'hcf7b8c;
		12'd0539: rd_data_1 <= 24'hc7848c;
		12'd0540: rd_data_1 <= 24'h9e787a;
		12'd0541: rd_data_1 <= 24'h807d7d;
		12'd0542: rd_data_1 <= 24'h56757a;
		12'd0543: rd_data_1 <= 24'h2e606b;
		12'd0544: rd_data_1 <= 24'h336c78;
		12'd0545: rd_data_1 <= 24'h275762;
		12'd0546: rd_data_1 <= 24'h133842;
		12'd0547: rd_data_1 <= 24'h27636b;
		12'd0548: rd_data_1 <= 24'h408f8e;
		12'd0549: rd_data_1 <= 24'h338e85;
		12'd0550: rd_data_1 <= 24'h3e958b;
		12'd0551: rd_data_1 <= 24'h39877d;
		12'd0552: rd_data_1 <= 24'h2d7c70;
		12'd0553: rd_data_1 <= 24'h36887b;
		12'd0554: rd_data_1 <= 24'h4b9a8f;
		12'd0555: rd_data_1 <= 24'h458f89;
		12'd0556: rd_data_1 <= 24'h37807d;
		12'd0557: rd_data_1 <= 24'h4e9297;
		12'd0558: rd_data_1 <= 24'h4e798a;
		12'd0559: rd_data_1 <= 24'h3d3f63;
		12'd0560: rd_data_1 <= 24'h3f0d51;
		12'd0561: rd_data_1 <= 24'h730977;
		12'd0562: rd_data_1 <= 24'h7f007e;
		12'd0563: rd_data_1 <= 24'h7e017d;
		12'd0564: rd_data_1 <= 24'h7e017d;
		12'd0565: rd_data_1 <= 24'h7e007e;
		12'd0566: rd_data_1 <= 24'h7e007e;
		12'd0567: rd_data_1 <= 24'h7e007e;
		12'd0568: rd_data_1 <= 24'h7e007e;
		12'd0569: rd_data_1 <= 24'h7e007e;
		12'd0570: rd_data_1 <= 24'h7e007e;
		12'd0571: rd_data_1 <= 24'h7e007e;
		12'd0572: rd_data_1 <= 24'h7e007e;
		12'd0573: rd_data_1 <= 24'h7f007f;
		12'd0574: rd_data_1 <= 24'h7f007f;
		12'd0575: rd_data_1 <= 24'h7f007f;
		12'd0576: rd_data_1 <= 24'h7f007f;
		12'd0577: rd_data_1 <= 24'h7f007f;
		12'd0578: rd_data_1 <= 24'h7f007f;
		12'd0579: rd_data_1 <= 24'h7f007f;
		12'd0580: rd_data_1 <= 24'h7f007f;
		12'd0581: rd_data_1 <= 24'h7f007f;
		12'd0582: rd_data_1 <= 24'h7f007f;
		12'd0583: rd_data_1 <= 24'h7f007f;
		12'd0584: rd_data_1 <= 24'h800080;
		12'd0585: rd_data_1 <= 24'h800080;
		12'd0586: rd_data_1 <= 24'h80007d;
		12'd0587: rd_data_1 <= 24'h80007e;
		12'd0588: rd_data_1 <= 24'h7c0080;
		12'd0589: rd_data_1 <= 24'h7d0080;
		12'd0590: rd_data_1 <= 24'h80007f;
		12'd0591: rd_data_1 <= 24'h82007d;
		12'd0592: rd_data_1 <= 24'h7e0378;
		12'd0593: rd_data_1 <= 24'h760977;
		12'd0594: rd_data_1 <= 24'h641478;
		12'd0595: rd_data_1 <= 24'h2d0550;
		12'd0596: rd_data_1 <= 24'h151936;
		12'd0597: rd_data_1 <= 24'h355655;
		12'd0598: rd_data_1 <= 24'h496960;
		12'd0599: rd_data_1 <= 24'h495f59;
		12'd0600: rd_data_1 <= 24'h4e585c;
		12'd0601: rd_data_1 <= 24'h4f555e;
		12'd0602: rd_data_1 <= 24'h535859;
		12'd0603: rd_data_1 <= 24'h565e55;
		12'd0604: rd_data_1 <= 24'h4f6251;
		12'd0605: rd_data_1 <= 24'h4b6754;
		12'd0606: rd_data_1 <= 24'h275148;
		12'd0607: rd_data_1 <= 24'h153f41;
		12'd0608: rd_data_1 <= 24'h123841;
		12'd0609: rd_data_1 <= 24'h2a606e;
		12'd0610: rd_data_1 <= 24'h4a98a1;
		12'd0611: rd_data_1 <= 24'h3a9294;
		12'd0612: rd_data_1 <= 24'h1f7a75;
		12'd0613: rd_data_1 <= 24'h1e746c;
		12'd0614: rd_data_1 <= 24'h47958f;
		12'd0615: rd_data_1 <= 24'h2e7269;
		12'd0616: rd_data_1 <= 24'h0e574b;
		12'd0617: rd_data_1 <= 24'h439d8f;
		12'd0618: rd_data_1 <= 24'h3e9087;
		12'd0619: rd_data_1 <= 24'h276c6b;
		12'd0620: rd_data_1 <= 24'h115356;
		12'd0621: rd_data_1 <= 24'h387b82;
		12'd0622: rd_data_1 <= 24'h528796;
		12'd0623: rd_data_1 <= 24'h576e8b;
		12'd0624: rd_data_1 <= 24'h210141;
		12'd0625: rd_data_1 <= 24'h700c78;
		12'd0626: rd_data_1 <= 24'h80007e;
		12'd0627: rd_data_1 <= 24'h7e017d;
		12'd0628: rd_data_1 <= 24'h7e017d;
		12'd0629: rd_data_1 <= 24'h7f007d;
		12'd0630: rd_data_1 <= 24'h7f007d;
		12'd0631: rd_data_1 <= 24'h7f007d;
		12'd0632: rd_data_1 <= 24'h7f007d;
		12'd0633: rd_data_1 <= 24'h7f007d;
		12'd0634: rd_data_1 <= 24'h7f007d;
		12'd0635: rd_data_1 <= 24'h7f007d;
		12'd0636: rd_data_1 <= 24'h7f007d;
		12'd0637: rd_data_1 <= 24'h7f007f;
		12'd0638: rd_data_1 <= 24'h7f007f;
		12'd0639: rd_data_1 <= 24'h7f007f;
		12'd0640: rd_data_1 <= 24'h7f007f;
		12'd0641: rd_data_1 <= 24'h7f007f;
		12'd0642: rd_data_1 <= 24'h7f007f;
		12'd0643: rd_data_1 <= 24'h7f007f;
		12'd0644: rd_data_1 <= 24'h7f007f;
		12'd0645: rd_data_1 <= 24'h7f007f;
		12'd0646: rd_data_1 <= 24'h7f007f;
		12'd0647: rd_data_1 <= 24'h7f007f;
		12'd0648: rd_data_1 <= 24'h7f007f;
		12'd0649: rd_data_1 <= 24'h7f007f;
		12'd0650: rd_data_1 <= 24'h7f007e;
		12'd0651: rd_data_1 <= 24'h7f007f;
		12'd0652: rd_data_1 <= 24'h7d007e;
		12'd0653: rd_data_1 <= 24'h7d007f;
		12'd0654: rd_data_1 <= 24'h80007e;
		12'd0655: rd_data_1 <= 24'h83007f;
		12'd0656: rd_data_1 <= 24'h7e0077;
		12'd0657: rd_data_1 <= 24'h7d017b;
		12'd0658: rd_data_1 <= 24'h6d0378;
		12'd0659: rd_data_1 <= 24'h692b85;
		12'd0660: rd_data_1 <= 24'h7c8caf;
		12'd0661: rd_data_1 <= 24'h366c65;
		12'd0662: rd_data_1 <= 24'h185641;
		12'd0663: rd_data_1 <= 24'h0f4633;
		12'd0664: rd_data_1 <= 24'h002b24;
		12'd0665: rd_data_1 <= 24'h073736;
		12'd0666: rd_data_1 <= 24'h14413a;
		12'd0667: rd_data_1 <= 24'h103c2c;
		12'd0668: rd_data_1 <= 24'h0d3f28;
		12'd0669: rd_data_1 <= 24'h093720;
		12'd0670: rd_data_1 <= 24'h306c5f;
		12'd0671: rd_data_1 <= 24'h46908e;
		12'd0672: rd_data_1 <= 24'h459497;
		12'd0673: rd_data_1 <= 24'h53a9ae;
		12'd0674: rd_data_1 <= 24'h3e989b;
		12'd0675: rd_data_1 <= 24'h359392;
		12'd0676: rd_data_1 <= 24'h257e7b;
		12'd0677: rd_data_1 <= 24'h1c6a66;
		12'd0678: rd_data_1 <= 24'h397976;
		12'd0679: rd_data_1 <= 24'h2a5856;
		12'd0680: rd_data_1 <= 24'h1e5e58;
		12'd0681: rd_data_1 <= 24'h3d9d93;
		12'd0682: rd_data_1 <= 24'h2c817c;
		12'd0683: rd_data_1 <= 24'h0c4d50;
		12'd0684: rd_data_1 <= 24'h114d52;
		12'd0685: rd_data_1 <= 24'h1a575e;
		12'd0686: rd_data_1 <= 24'h548893;
		12'd0687: rd_data_1 <= 24'h4f6e83;
		12'd0688: rd_data_1 <= 24'h1d053d;
		12'd0689: rd_data_1 <= 24'h700c78;
		12'd0690: rd_data_1 <= 24'h80007e;
		12'd0691: rd_data_1 <= 24'h7e017d;
		12'd0692: rd_data_1 <= 24'h7e017d;
		12'd0693: rd_data_1 <= 24'h7f007d;
		12'd0694: rd_data_1 <= 24'h7f007d;
		12'd0695: rd_data_1 <= 24'h7f007d;
		12'd0696: rd_data_1 <= 24'h7f007d;
		12'd0697: rd_data_1 <= 24'h7f007d;
		12'd0698: rd_data_1 <= 24'h7f007d;
		12'd0699: rd_data_1 <= 24'h7f007d;
		12'd0700: rd_data_1 <= 24'h7f007d;
		12'd0701: rd_data_1 <= 24'h7f007f;
		12'd0702: rd_data_1 <= 24'h7f007f;
		12'd0703: rd_data_1 <= 24'h7f007f;
		12'd0704: rd_data_1 <= 24'h7f007f;
		12'd0705: rd_data_1 <= 24'h7f007f;
		12'd0706: rd_data_1 <= 24'h7f007f;
		12'd0707: rd_data_1 <= 24'h7f007f;
		12'd0708: rd_data_1 <= 24'h7f007f;
		12'd0709: rd_data_1 <= 24'h7f007f;
		12'd0710: rd_data_1 <= 24'h7f007f;
		12'd0711: rd_data_1 <= 24'h7f007f;
		12'd0712: rd_data_1 <= 24'h7f007f;
		12'd0713: rd_data_1 <= 24'h7f007f;
		12'd0714: rd_data_1 <= 24'h7f007f;
		12'd0715: rd_data_1 <= 24'h7f007f;
		12'd0716: rd_data_1 <= 24'h7d007e;
		12'd0717: rd_data_1 <= 24'h7d007e;
		12'd0718: rd_data_1 <= 24'h80007e;
		12'd0719: rd_data_1 <= 24'h82007e;
		12'd0720: rd_data_1 <= 24'h870382;
		12'd0721: rd_data_1 <= 24'h790077;
		12'd0722: rd_data_1 <= 24'h740379;
		12'd0723: rd_data_1 <= 24'h7e3793;
		12'd0724: rd_data_1 <= 24'h7f91b3;
		12'd0725: rd_data_1 <= 24'h65bcb1;
		12'd0726: rd_data_1 <= 24'h6cd5bf;
		12'd0727: rd_data_1 <= 24'h60c2af;
		12'd0728: rd_data_1 <= 24'h2a7a71;
		12'd0729: rd_data_1 <= 24'h327270;
		12'd0730: rd_data_1 <= 24'h427d74;
		12'd0731: rd_data_1 <= 24'h4c8d7d;
		12'd0732: rd_data_1 <= 24'h54a190;
		12'd0733: rd_data_1 <= 24'h489e90;
		12'd0734: rd_data_1 <= 24'h3d8b85;
		12'd0735: rd_data_1 <= 24'h1c6664;
		12'd0736: rd_data_1 <= 24'h32908a;
		12'd0737: rd_data_1 <= 24'h68d8d1;
		12'd0738: rd_data_1 <= 24'h59c3be;
		12'd0739: rd_data_1 <= 24'h3e9c98;
		12'd0740: rd_data_1 <= 24'h419291;
		12'd0741: rd_data_1 <= 24'h347b7b;
		12'd0742: rd_data_1 <= 24'h002c30;
		12'd0743: rd_data_1 <= 24'h1a363e;
		12'd0744: rd_data_1 <= 24'h569c9f;
		12'd0745: rd_data_1 <= 24'h3b9b96;
		12'd0746: rd_data_1 <= 24'h247c7a;
		12'd0747: rd_data_1 <= 24'h0b4b50;
		12'd0748: rd_data_1 <= 24'h0d444c;
		12'd0749: rd_data_1 <= 24'h225b61;
		12'd0750: rd_data_1 <= 24'h5f8e96;
		12'd0751: rd_data_1 <= 24'h4d6676;
		12'd0752: rd_data_1 <= 24'h1a0132;
		12'd0753: rd_data_1 <= 24'h710d77;
		12'd0754: rd_data_1 <= 24'h80007e;
		12'd0755: rd_data_1 <= 24'h7e017d;
		12'd0756: rd_data_1 <= 24'h7e017d;
		12'd0757: rd_data_1 <= 24'h7f007d;
		12'd0758: rd_data_1 <= 24'h7f007d;
		12'd0759: rd_data_1 <= 24'h7f007d;
		12'd0760: rd_data_1 <= 24'h7f007d;
		12'd0761: rd_data_1 <= 24'h7f007d;
		12'd0762: rd_data_1 <= 24'h7f007d;
		12'd0763: rd_data_1 <= 24'h7f007d;
		12'd0764: rd_data_1 <= 24'h7f007d;
		12'd0765: rd_data_1 <= 24'h7f007f;
		12'd0766: rd_data_1 <= 24'h7f007f;
		12'd0767: rd_data_1 <= 24'h7f007f;
		12'd0768: rd_data_1 <= 24'h7f007f;
		12'd0769: rd_data_1 <= 24'h7f007f;
		12'd0770: rd_data_1 <= 24'h7f007f;
		12'd0771: rd_data_1 <= 24'h7f007f;
		12'd0772: rd_data_1 <= 24'h7f007f;
		12'd0773: rd_data_1 <= 24'h7f007f;
		12'd0774: rd_data_1 <= 24'h7f007f;
		12'd0775: rd_data_1 <= 24'h7f007f;
		12'd0776: rd_data_1 <= 24'h7f007f;
		12'd0777: rd_data_1 <= 24'h7f007f;
		12'd0778: rd_data_1 <= 24'h7f007f;
		12'd0779: rd_data_1 <= 24'h7f007f;
		12'd0780: rd_data_1 <= 24'h7d007e;
		12'd0781: rd_data_1 <= 24'h7e007e;
		12'd0782: rd_data_1 <= 24'h80007e;
		12'd0783: rd_data_1 <= 24'h81007d;
		12'd0784: rd_data_1 <= 24'h880684;
		12'd0785: rd_data_1 <= 24'h7e027c;
		12'd0786: rd_data_1 <= 24'h7e037e;
		12'd0787: rd_data_1 <= 24'h5f0c6c;
		12'd0788: rd_data_1 <= 24'h404c71;
		12'd0789: rd_data_1 <= 24'h2d827a;
		12'd0790: rd_data_1 <= 24'h52bba5;
		12'd0791: rd_data_1 <= 24'h6fd5c0;
		12'd0792: rd_data_1 <= 24'h52a89e;
		12'd0793: rd_data_1 <= 24'h256d6c;
		12'd0794: rd_data_1 <= 24'h134742;
		12'd0795: rd_data_1 <= 24'h26574f;
		12'd0796: rd_data_1 <= 24'h3c696e;
		12'd0797: rd_data_1 <= 24'h3d6775;
		12'd0798: rd_data_1 <= 24'h164f56;
		12'd0799: rd_data_1 <= 24'h24716c;
		12'd0800: rd_data_1 <= 24'h3d9b92;
		12'd0801: rd_data_1 <= 24'h3ea69c;
		12'd0802: rd_data_1 <= 24'h68cfc6;
		12'd0803: rd_data_1 <= 24'h5dbcb6;
		12'd0804: rd_data_1 <= 24'h3b8c8b;
		12'd0805: rd_data_1 <= 24'h327377;
		12'd0806: rd_data_1 <= 24'h08313c;
		12'd0807: rd_data_1 <= 24'h223d4d;
		12'd0808: rd_data_1 <= 24'h63979f;
		12'd0809: rd_data_1 <= 24'h439c99;
		12'd0810: rd_data_1 <= 24'h338e8b;
		12'd0811: rd_data_1 <= 24'h135e5f;
		12'd0812: rd_data_1 <= 24'h0a4d52;
		12'd0813: rd_data_1 <= 24'h337176;
		12'd0814: rd_data_1 <= 24'h57838e;
		12'd0815: rd_data_1 <= 24'h424a61;
		12'd0816: rd_data_1 <= 24'h350a45;
		12'd0817: rd_data_1 <= 24'h720b75;
		12'd0818: rd_data_1 <= 24'h7f007e;
		12'd0819: rd_data_1 <= 24'h7e017d;
		12'd0820: rd_data_1 <= 24'h7e017d;
		12'd0821: rd_data_1 <= 24'h7f007d;
		12'd0822: rd_data_1 <= 24'h7f007d;
		12'd0823: rd_data_1 <= 24'h7f007d;
		12'd0824: rd_data_1 <= 24'h7f007d;
		12'd0825: rd_data_1 <= 24'h7f007d;
		12'd0826: rd_data_1 <= 24'h7f007d;
		12'd0827: rd_data_1 <= 24'h7f007d;
		12'd0828: rd_data_1 <= 24'h7f007d;
		12'd0829: rd_data_1 <= 24'h7f007f;
		12'd0830: rd_data_1 <= 24'h7f007f;
		12'd0831: rd_data_1 <= 24'h7f007f;
		12'd0832: rd_data_1 <= 24'h7f007f;
		12'd0833: rd_data_1 <= 24'h7f007f;
		12'd0834: rd_data_1 <= 24'h7f007f;
		12'd0835: rd_data_1 <= 24'h7f007f;
		12'd0836: rd_data_1 <= 24'h7f007f;
		12'd0837: rd_data_1 <= 24'h7f007f;
		12'd0838: rd_data_1 <= 24'h7f007f;
		12'd0839: rd_data_1 <= 24'h7f007f;
		12'd0840: rd_data_1 <= 24'h7f007f;
		12'd0841: rd_data_1 <= 24'h7f007f;
		12'd0842: rd_data_1 <= 24'h7f007f;
		12'd0843: rd_data_1 <= 24'h7f007f;
		12'd0844: rd_data_1 <= 24'h7e007f;
		12'd0845: rd_data_1 <= 24'h7f007f;
		12'd0846: rd_data_1 <= 24'h81007f;
		12'd0847: rd_data_1 <= 24'h83007f;
		12'd0848: rd_data_1 <= 24'h83007d;
		12'd0849: rd_data_1 <= 24'h80007d;
		12'd0850: rd_data_1 <= 24'h82017e;
		12'd0851: rd_data_1 <= 24'h680a6e;
		12'd0852: rd_data_1 <= 24'h53517b;
		12'd0853: rd_data_1 <= 24'h4b9490;
		12'd0854: rd_data_1 <= 24'h5cbdaa;
		12'd0855: rd_data_1 <= 24'h6ed2be;
		12'd0856: rd_data_1 <= 24'h5ab4ab;
		12'd0857: rd_data_1 <= 24'h4c9696;
		12'd0858: rd_data_1 <= 24'h669d9d;
		12'd0859: rd_data_1 <= 24'h2c474e;
		12'd0860: rd_data_1 <= 24'h110327;
		12'd0861: rd_data_1 <= 24'h1d0337;
		12'd0862: rd_data_1 <= 24'h1c344d;
		12'd0863: rd_data_1 <= 24'h3d8c84;
		12'd0864: rd_data_1 <= 24'h459d91;
		12'd0865: rd_data_1 <= 24'h33867e;
		12'd0866: rd_data_1 <= 24'h52aea4;
		12'd0867: rd_data_1 <= 24'h5dbfb5;
		12'd0868: rd_data_1 <= 24'h3f908f;
		12'd0869: rd_data_1 <= 24'h346c76;
		12'd0870: rd_data_1 <= 24'h132e41;
		12'd0871: rd_data_1 <= 24'h252f48;
		12'd0872: rd_data_1 <= 24'h4f6f7d;
		12'd0873: rd_data_1 <= 24'h3f8787;
		12'd0874: rd_data_1 <= 24'h419891;
		12'd0875: rd_data_1 <= 24'h2e807c;
		12'd0876: rd_data_1 <= 24'h217170;
		12'd0877: rd_data_1 <= 24'h4c8f95;
		12'd0878: rd_data_1 <= 24'h46677c;
		12'd0879: rd_data_1 <= 24'h13022a;
		12'd0880: rd_data_1 <= 24'h55135c;
		12'd0881: rd_data_1 <= 24'h760776;
		12'd0882: rd_data_1 <= 24'h80007e;
		12'd0883: rd_data_1 <= 24'h7f007d;
		12'd0884: rd_data_1 <= 24'h7f007d;
		12'd0885: rd_data_1 <= 24'h7f007d;
		12'd0886: rd_data_1 <= 24'h7f007d;
		12'd0887: rd_data_1 <= 24'h7f007d;
		12'd0888: rd_data_1 <= 24'h7f007d;
		12'd0889: rd_data_1 <= 24'h7f007d;
		12'd0890: rd_data_1 <= 24'h7f007d;
		12'd0891: rd_data_1 <= 24'h7f007d;
		12'd0892: rd_data_1 <= 24'h7f007d;
		12'd0893: rd_data_1 <= 24'h7f007f;
		12'd0894: rd_data_1 <= 24'h7f007f;
		12'd0895: rd_data_1 <= 24'h7f007f;
		12'd0896: rd_data_1 <= 24'h7f007f;
		12'd0897: rd_data_1 <= 24'h7f007f;
		12'd0898: rd_data_1 <= 24'h7f007f;
		12'd0899: rd_data_1 <= 24'h7f007f;
		12'd0900: rd_data_1 <= 24'h7f007f;
		12'd0901: rd_data_1 <= 24'h7f007f;
		12'd0902: rd_data_1 <= 24'h7f007f;
		12'd0903: rd_data_1 <= 24'h7f007f;
		12'd0904: rd_data_1 <= 24'h7f007f;
		12'd0905: rd_data_1 <= 24'h7f007f;
		12'd0906: rd_data_1 <= 24'h7f007f;
		12'd0907: rd_data_1 <= 24'h7f007f;
		12'd0908: rd_data_1 <= 24'h7e007f;
		12'd0909: rd_data_1 <= 24'h7f007f;
		12'd0910: rd_data_1 <= 24'h81007f;
		12'd0911: rd_data_1 <= 24'h83007f;
		12'd0912: rd_data_1 <= 24'h84007e;
		12'd0913: rd_data_1 <= 24'h83007e;
		12'd0914: rd_data_1 <= 24'h83007e;
		12'd0915: rd_data_1 <= 24'h6d086e;
		12'd0916: rd_data_1 <= 24'h604b7b;
		12'd0917: rd_data_1 <= 24'h729fa5;
		12'd0918: rd_data_1 <= 24'h7cc8bc;
		12'd0919: rd_data_1 <= 24'h6ac4b4;
		12'd0920: rd_data_1 <= 24'h78d6cd;
		12'd0921: rd_data_1 <= 24'h58aaab;
		12'd0922: rd_data_1 <= 24'h59898f;
		12'd0923: rd_data_1 <= 24'h34384c;
		12'd0924: rd_data_1 <= 24'h390b42;
		12'd0925: rd_data_1 <= 24'h541963;
		12'd0926: rd_data_1 <= 24'h51597c;
		12'd0927: rd_data_1 <= 24'h6ab9b0;
		12'd0928: rd_data_1 <= 24'h62bbaa;
		12'd0929: rd_data_1 <= 24'h4a998e;
		12'd0930: rd_data_1 <= 24'h59b6aa;
		12'd0931: rd_data_1 <= 24'h52b5a9;
		12'd0932: rd_data_1 <= 24'h3d7f83;
		12'd0933: rd_data_1 <= 24'h445a71;
		12'd0934: rd_data_1 <= 24'h3c3459;
		12'd0935: rd_data_1 <= 24'h2a193f;
		12'd0936: rd_data_1 <= 24'h283042;
		12'd0937: rd_data_1 <= 24'h578681;
		12'd0938: rd_data_1 <= 24'h478479;
		12'd0939: rd_data_1 <= 24'h4d8885;
		12'd0940: rd_data_1 <= 24'h4b8086;
		12'd0941: rd_data_1 <= 24'h5a8194;
		12'd0942: rd_data_1 <= 24'h55537c;
		12'd0943: rd_data_1 <= 24'h380142;
		12'd0944: rd_data_1 <= 24'h680a66;
		12'd0945: rd_data_1 <= 24'h7b0479;
		12'd0946: rd_data_1 <= 24'h80007e;
		12'd0947: rd_data_1 <= 24'h7f007d;
		12'd0948: rd_data_1 <= 24'h7f007d;
		12'd0949: rd_data_1 <= 24'h7f007d;
		12'd0950: rd_data_1 <= 24'h7f007d;
		12'd0951: rd_data_1 <= 24'h7f007d;
		12'd0952: rd_data_1 <= 24'h7f007d;
		12'd0953: rd_data_1 <= 24'h7f007d;
		12'd0954: rd_data_1 <= 24'h7f007d;
		12'd0955: rd_data_1 <= 24'h7f007d;
		12'd0956: rd_data_1 <= 24'h7f007d;
		12'd0957: rd_data_1 <= 24'h7f007f;
		12'd0958: rd_data_1 <= 24'h7f007f;
		12'd0959: rd_data_1 <= 24'h7f007f;
		12'd0960: rd_data_1 <= 24'h7f007f;
		12'd0961: rd_data_1 <= 24'h7f007f;
		12'd0962: rd_data_1 <= 24'h7f007f;
		12'd0963: rd_data_1 <= 24'h7f007f;
		12'd0964: rd_data_1 <= 24'h7f007f;
		12'd0965: rd_data_1 <= 24'h7f007f;
		12'd0966: rd_data_1 <= 24'h7f007f;
		12'd0967: rd_data_1 <= 24'h7f007f;
		12'd0968: rd_data_1 <= 24'h7f007f;
		12'd0969: rd_data_1 <= 24'h7f007f;
		12'd0970: rd_data_1 <= 24'h7f007f;
		12'd0971: rd_data_1 <= 24'h7f007f;
		12'd0972: rd_data_1 <= 24'h7e007f;
		12'd0973: rd_data_1 <= 24'h7f007f;
		12'd0974: rd_data_1 <= 24'h81007f;
		12'd0975: rd_data_1 <= 24'h83007f;
		12'd0976: rd_data_1 <= 24'h85007f;
		12'd0977: rd_data_1 <= 24'h84007e;
		12'd0978: rd_data_1 <= 24'h83007e;
		12'd0979: rd_data_1 <= 24'h730b73;
		12'd0980: rd_data_1 <= 24'h481a54;
		12'd0981: rd_data_1 <= 24'h606978;
		12'd0982: rd_data_1 <= 24'h7ba6a5;
		12'd0983: rd_data_1 <= 24'h6fb1a9;
		12'd0984: rd_data_1 <= 24'h5db5ae;
		12'd0985: rd_data_1 <= 24'h50a2a5;
		12'd0986: rd_data_1 <= 24'h527683;
		12'd0987: rd_data_1 <= 24'h362544;
		12'd0988: rd_data_1 <= 24'h48084e;
		12'd0989: rd_data_1 <= 24'h59146c;
		12'd0990: rd_data_1 <= 24'h40416c;
		12'd0991: rd_data_1 <= 24'h5ba89f;
		12'd0992: rd_data_1 <= 24'h71cbb7;
		12'd0993: rd_data_1 <= 24'h74c7b6;
		12'd0994: rd_data_1 <= 24'h70cdbd;
		12'd0995: rd_data_1 <= 24'h56afa6;
		12'd0996: rd_data_1 <= 24'h305463;
		12'd0997: rd_data_1 <= 24'h230631;
		12'd0998: rd_data_1 <= 24'h59235c;
		12'd0999: rd_data_1 <= 24'h4e1e55;
		12'd1000: rd_data_1 <= 24'h6d5873;
		12'd1001: rd_data_1 <= 24'h77837d;
		12'd1002: rd_data_1 <= 24'h40534b;
		12'd1003: rd_data_1 <= 24'h879198;
		12'd1004: rd_data_1 <= 24'h44455e;
		12'd1005: rd_data_1 <= 24'h9f8ebc;
		12'd1006: rd_data_1 <= 24'h481258;
		12'd1007: rd_data_1 <= 24'h6d0769;
		12'd1008: rd_data_1 <= 24'h7b0072;
		12'd1009: rd_data_1 <= 24'h7e017b;
		12'd1010: rd_data_1 <= 24'h7f007d;
		12'd1011: rd_data_1 <= 24'h7f007d;
		12'd1012: rd_data_1 <= 24'h7f007d;
		12'd1013: rd_data_1 <= 24'h7f007d;
		12'd1014: rd_data_1 <= 24'h7f007d;
		12'd1015: rd_data_1 <= 24'h7f007d;
		12'd1016: rd_data_1 <= 24'h7f007d;
		12'd1017: rd_data_1 <= 24'h7f007d;
		12'd1018: rd_data_1 <= 24'h7f007d;
		12'd1019: rd_data_1 <= 24'h7f007d;
		12'd1020: rd_data_1 <= 24'h7f007d;
		12'd1021: rd_data_1 <= 24'h7f007f;
		12'd1022: rd_data_1 <= 24'h7f007f;
		12'd1023: rd_data_1 <= 24'h7f007f;
		12'd1024: rd_data_1 <= 24'h7f007f;
		12'd1025: rd_data_1 <= 24'h7f007f;
		12'd1026: rd_data_1 <= 24'h7f007f;
		12'd1027: rd_data_1 <= 24'h7f007f;
		12'd1028: rd_data_1 <= 24'h7f007f;
		12'd1029: rd_data_1 <= 24'h7f007f;
		12'd1030: rd_data_1 <= 24'h7f007f;
		12'd1031: rd_data_1 <= 24'h7f007f;
		12'd1032: rd_data_1 <= 24'h7f007f;
		12'd1033: rd_data_1 <= 24'h7f007f;
		12'd1034: rd_data_1 <= 24'h7f007f;
		12'd1035: rd_data_1 <= 24'h7f007f;
		12'd1036: rd_data_1 <= 24'h7e007f;
		12'd1037: rd_data_1 <= 24'h7f007f;
		12'd1038: rd_data_1 <= 24'h81007f;
		12'd1039: rd_data_1 <= 24'h83007f;
		12'd1040: rd_data_1 <= 24'h850083;
		12'd1041: rd_data_1 <= 24'h850083;
		12'd1042: rd_data_1 <= 24'h83017f;
		12'd1043: rd_data_1 <= 24'h760875;
		12'd1044: rd_data_1 <= 24'h55115b;
		12'd1045: rd_data_1 <= 24'hc6abc6;
		12'd1046: rd_data_1 <= 24'h565a69;
		12'd1047: rd_data_1 <= 24'h94a1ab;
		12'd1048: rd_data_1 <= 24'h51737e;
		12'd1049: rd_data_1 <= 24'h315569;
		12'd1050: rd_data_1 <= 24'h352e52;
		12'd1051: rd_data_1 <= 24'h410c4a;
		12'd1052: rd_data_1 <= 24'h681671;
		12'd1053: rd_data_1 <= 24'h5b1273;
		12'd1054: rd_data_1 <= 24'h4e4473;
		12'd1055: rd_data_1 <= 24'h5e9494;
		12'd1056: rd_data_1 <= 24'h6faea4;
		12'd1057: rd_data_1 <= 24'h74a9a0;
		12'd1058: rd_data_1 <= 24'h76ada7;
		12'd1059: rd_data_1 <= 24'h68939b;
		12'd1060: rd_data_1 <= 24'h423d60;
		12'd1061: rd_data_1 <= 24'h410343;
		12'd1062: rd_data_1 <= 24'h691165;
		12'd1063: rd_data_1 <= 24'h620c63;
		12'd1064: rd_data_1 <= 24'h490647;
		12'd1065: rd_data_1 <= 24'h24001f;
		12'd1066: rd_data_1 <= 24'h280225;
		12'd1067: rd_data_1 <= 24'h29002b;
		12'd1068: rd_data_1 <= 24'h31003a;
		12'd1069: rd_data_1 <= 24'h3c0048;
		12'd1070: rd_data_1 <= 24'h6b1070;
		12'd1071: rd_data_1 <= 24'h800577;
		12'd1072: rd_data_1 <= 24'h86027c;
		12'd1073: rd_data_1 <= 24'h80007b;
		12'd1074: rd_data_1 <= 24'h7f007d;
		12'd1075: rd_data_1 <= 24'h7f007d;
		12'd1076: rd_data_1 <= 24'h7f007d;
		12'd1077: rd_data_1 <= 24'h7f007d;
		12'd1078: rd_data_1 <= 24'h7f007d;
		12'd1079: rd_data_1 <= 24'h7f007d;
		12'd1080: rd_data_1 <= 24'h7f007d;
		12'd1081: rd_data_1 <= 24'h7f007d;
		12'd1082: rd_data_1 <= 24'h7f007d;
		12'd1083: rd_data_1 <= 24'h7f007d;
		12'd1084: rd_data_1 <= 24'h7f007d;
		12'd1085: rd_data_1 <= 24'h7f007f;
		12'd1086: rd_data_1 <= 24'h7f007f;
		12'd1087: rd_data_1 <= 24'h7f007f;
		12'd1088: rd_data_1 <= 24'h7f007f;
		12'd1089: rd_data_1 <= 24'h7f007f;
		12'd1090: rd_data_1 <= 24'h7f007f;
		12'd1091: rd_data_1 <= 24'h7f007f;
		12'd1092: rd_data_1 <= 24'h7f007f;
		12'd1093: rd_data_1 <= 24'h7f007f;
		12'd1094: rd_data_1 <= 24'h7f007f;
		12'd1095: rd_data_1 <= 24'h7f007f;
		12'd1096: rd_data_1 <= 24'h7f007f;
		12'd1097: rd_data_1 <= 24'h7f007f;
		12'd1098: rd_data_1 <= 24'h7f007f;
		12'd1099: rd_data_1 <= 24'h7f007f;
		12'd1100: rd_data_1 <= 24'h7e007f;
		12'd1101: rd_data_1 <= 24'h7f007f;
		12'd1102: rd_data_1 <= 24'h81007f;
		12'd1103: rd_data_1 <= 24'h830080;
		12'd1104: rd_data_1 <= 24'h850087;
		12'd1105: rd_data_1 <= 24'h85008a;
		12'd1106: rd_data_1 <= 24'h810183;
		12'd1107: rd_data_1 <= 24'h77077b;
		12'd1108: rd_data_1 <= 24'h6b106d;
		12'd1109: rd_data_1 <= 24'h3c0040;
		12'd1110: rd_data_1 <= 24'h240029;
		12'd1111: rd_data_1 <= 24'h1f0025;
		12'd1112: rd_data_1 <= 24'h1f0027;
		12'd1113: rd_data_1 <= 24'h26002f;
		12'd1114: rd_data_1 <= 24'h520d59;
		12'd1115: rd_data_1 <= 24'h6f1177;
		12'd1116: rd_data_1 <= 24'h6a0979;
		12'd1117: rd_data_1 <= 24'h570a71;
		12'd1118: rd_data_1 <= 24'had8ebe;
		12'd1119: rd_data_1 <= 24'h76818e;
		12'd1120: rd_data_1 <= 24'h75818d;
		12'd1121: rd_data_1 <= 24'h878691;
		12'd1122: rd_data_1 <= 24'h797283;
		12'd1123: rd_data_1 <= 24'h9980a2;
		12'd1124: rd_data_1 <= 24'h34003f;
		12'd1125: rd_data_1 <= 24'h6c116e;
		12'd1126: rd_data_1 <= 24'h750575;
		12'd1127: rd_data_1 <= 24'h7b027b;
		12'd1128: rd_data_1 <= 24'h790479;
		12'd1129: rd_data_1 <= 24'h740a73;
		12'd1130: rd_data_1 <= 24'h730b72;
		12'd1131: rd_data_1 <= 24'h740975;
		12'd1132: rd_data_1 <= 24'h750978;
		12'd1133: rd_data_1 <= 24'h75077a;
		12'd1134: rd_data_1 <= 24'h780379;
		12'd1135: rd_data_1 <= 24'h7d007c;
		12'd1136: rd_data_1 <= 24'h7f007c;
		12'd1137: rd_data_1 <= 24'h7f007d;
		12'd1138: rd_data_1 <= 24'h7f007f;
		12'd1139: rd_data_1 <= 24'h7f007f;
		12'd1140: rd_data_1 <= 24'h7f007f;
		12'd1141: rd_data_1 <= 24'h7f007f;
		12'd1142: rd_data_1 <= 24'h7f007f;
		12'd1143: rd_data_1 <= 24'h7f007f;
		12'd1144: rd_data_1 <= 24'h7f007f;
		12'd1145: rd_data_1 <= 24'h7f007f;
		12'd1146: rd_data_1 <= 24'h7f007f;
		12'd1147: rd_data_1 <= 24'h7f007f;
		12'd1148: rd_data_1 <= 24'h7f007f;
		12'd1149: rd_data_1 <= 24'h7f007f;
		12'd1150: rd_data_1 <= 24'h7f007f;
		12'd1151: rd_data_1 <= 24'h7f007f;
		12'd1152: rd_data_1 <= 24'h7f007f;
		12'd1153: rd_data_1 <= 24'h7f007f;
		12'd1154: rd_data_1 <= 24'h7f007f;
		12'd1155: rd_data_1 <= 24'h7f007f;
		12'd1156: rd_data_1 <= 24'h7f007f;
		12'd1157: rd_data_1 <= 24'h7f007f;
		12'd1158: rd_data_1 <= 24'h7f007f;
		12'd1159: rd_data_1 <= 24'h7f007f;
		12'd1160: rd_data_1 <= 24'h7f007f;
		12'd1161: rd_data_1 <= 24'h7f007f;
		12'd1162: rd_data_1 <= 24'h7f007f;
		12'd1163: rd_data_1 <= 24'h7f007f;
		12'd1164: rd_data_1 <= 24'h7e007f;
		12'd1165: rd_data_1 <= 24'h7f007f;
		12'd1166: rd_data_1 <= 24'h81007f;
		12'd1167: rd_data_1 <= 24'h830080;
		12'd1168: rd_data_1 <= 24'h850086;
		12'd1169: rd_data_1 <= 24'h850088;
		12'd1170: rd_data_1 <= 24'h810182;
		12'd1171: rd_data_1 <= 24'h7a057b;
		12'd1172: rd_data_1 <= 24'h740a72;
		12'd1173: rd_data_1 <= 24'h6e0e6a;
		12'd1174: rd_data_1 <= 24'h681062;
		12'd1175: rd_data_1 <= 24'h66135d;
		12'd1176: rd_data_1 <= 24'h69125e;
		12'd1177: rd_data_1 <= 24'h6d0d64;
		12'd1178: rd_data_1 <= 24'h760875;
		12'd1179: rd_data_1 <= 24'h790581;
		12'd1180: rd_data_1 <= 24'h710583;
		12'd1181: rd_data_1 <= 24'h6a0d80;
		12'd1182: rd_data_1 <= 24'h41005b;
		12'd1183: rd_data_1 <= 24'h27003e;
		12'd1184: rd_data_1 <= 24'h240033;
		12'd1185: rd_data_1 <= 24'h2a0030;
		12'd1186: rd_data_1 <= 24'h330036;
		12'd1187: rd_data_1 <= 24'h49004c;
		12'd1188: rd_data_1 <= 24'h6e1170;
		12'd1189: rd_data_1 <= 24'h740574;
		12'd1190: rd_data_1 <= 24'h7d007d;
		12'd1191: rd_data_1 <= 24'h820081;
		12'd1192: rd_data_1 <= 24'h820082;
		12'd1193: rd_data_1 <= 24'h800080;
		12'd1194: rd_data_1 <= 24'h7f007f;
		12'd1195: rd_data_1 <= 24'h7f007f;
		12'd1196: rd_data_1 <= 24'h7f007f;
		12'd1197: rd_data_1 <= 24'h7f007f;
		12'd1198: rd_data_1 <= 24'h7f007e;
		12'd1199: rd_data_1 <= 24'h7e007e;
		12'd1200: rd_data_1 <= 24'h7e007e;
		12'd1201: rd_data_1 <= 24'h7f007f;
		12'd1202: rd_data_1 <= 24'h7f007f;
		12'd1203: rd_data_1 <= 24'h7f007f;
		12'd1204: rd_data_1 <= 24'h7f007f;
		12'd1205: rd_data_1 <= 24'h7f007f;
		12'd1206: rd_data_1 <= 24'h7f007f;
		12'd1207: rd_data_1 <= 24'h7f007f;
		12'd1208: rd_data_1 <= 24'h7f007f;
		12'd1209: rd_data_1 <= 24'h7f007f;
		12'd1210: rd_data_1 <= 24'h7f007f;
		12'd1211: rd_data_1 <= 24'h7f007f;
		12'd1212: rd_data_1 <= 24'h7f007f;
		12'd1213: rd_data_1 <= 24'h7f007f;
		12'd1214: rd_data_1 <= 24'h7f007f;
		12'd1215: rd_data_1 <= 24'h7f007f;
		12'd1216: rd_data_1 <= 24'h7f007f;
		12'd1217: rd_data_1 <= 24'h7f007f;
		12'd1218: rd_data_1 <= 24'h7f007f;
		12'd1219: rd_data_1 <= 24'h7f007f;
		12'd1220: rd_data_1 <= 24'h7f007f;
		12'd1221: rd_data_1 <= 24'h7f007f;
		12'd1222: rd_data_1 <= 24'h7f007f;
		12'd1223: rd_data_1 <= 24'h7f007f;
		12'd1224: rd_data_1 <= 24'h7f007f;
		12'd1225: rd_data_1 <= 24'h7f007f;
		12'd1226: rd_data_1 <= 24'h7f007f;
		12'd1227: rd_data_1 <= 24'h7f007f;
		12'd1228: rd_data_1 <= 24'h7e007f;
		12'd1229: rd_data_1 <= 24'h7f007f;
		12'd1230: rd_data_1 <= 24'h81007f;
		12'd1231: rd_data_1 <= 24'h81007f;
		12'd1232: rd_data_1 <= 24'h83007f;
		12'd1233: rd_data_1 <= 24'h84007f;
		12'd1234: rd_data_1 <= 24'h82017c;
		12'd1235: rd_data_1 <= 24'h80047a;
		12'd1236: rd_data_1 <= 24'h780373;
		12'd1237: rd_data_1 <= 24'h780672;
		12'd1238: rd_data_1 <= 24'h790b71;
		12'd1239: rd_data_1 <= 24'h780a70;
		12'd1240: rd_data_1 <= 24'h7d0776;
		12'd1241: rd_data_1 <= 24'h840781;
		12'd1242: rd_data_1 <= 24'h7f0283;
		12'd1243: rd_data_1 <= 24'h7c0186;
		12'd1244: rd_data_1 <= 24'h770086;
		12'd1245: rd_data_1 <= 24'h740284;
		12'd1246: rd_data_1 <= 24'h760883;
		12'd1247: rd_data_1 <= 24'h770e7f;
		12'd1248: rd_data_1 <= 24'h780e7e;
		12'd1249: rd_data_1 <= 24'h770a7d;
		12'd1250: rd_data_1 <= 24'h76077d;
		12'd1251: rd_data_1 <= 24'h76047a;
		12'd1252: rd_data_1 <= 24'h78037b;
		12'd1253: rd_data_1 <= 24'h7a017c;
		12'd1254: rd_data_1 <= 24'h7c007d;
		12'd1255: rd_data_1 <= 24'h7e007e;
		12'd1256: rd_data_1 <= 24'h7e007d;
		12'd1257: rd_data_1 <= 24'h7e007d;
		12'd1258: rd_data_1 <= 24'h7e007c;
		12'd1259: rd_data_1 <= 24'h7e007e;
		12'd1260: rd_data_1 <= 24'h7e007e;
		12'd1261: rd_data_1 <= 24'h7e007e;
		12'd1262: rd_data_1 <= 24'h7e007e;
		12'd1263: rd_data_1 <= 24'h7e007e;
		12'd1264: rd_data_1 <= 24'h7e007e;
		12'd1265: rd_data_1 <= 24'h7f007f;
		12'd1266: rd_data_1 <= 24'h7f007f;
		12'd1267: rd_data_1 <= 24'h7f007f;
		12'd1268: rd_data_1 <= 24'h7f007f;
		12'd1269: rd_data_1 <= 24'h7f007f;
		12'd1270: rd_data_1 <= 24'h7f007f;
		12'd1271: rd_data_1 <= 24'h7f007f;
		12'd1272: rd_data_1 <= 24'h7f007f;
		12'd1273: rd_data_1 <= 24'h7f007f;
		12'd1274: rd_data_1 <= 24'h7f007f;
		12'd1275: rd_data_1 <= 24'h7f007f;
		12'd1276: rd_data_1 <= 24'h7f007f;
		12'd1277: rd_data_1 <= 24'h7f007f;
		12'd1278: rd_data_1 <= 24'h7f007f;
		12'd1279: rd_data_1 <= 24'h7f007f;
		12'd1280: rd_data_1 <= 24'h7f007f;
		12'd1281: rd_data_1 <= 24'h7f007f;
		12'd1282: rd_data_1 <= 24'h7f007f;
		12'd1283: rd_data_1 <= 24'h7f007f;
		12'd1284: rd_data_1 <= 24'h7f007f;
		12'd1285: rd_data_1 <= 24'h7f007f;
		12'd1286: rd_data_1 <= 24'h7f007f;
		12'd1287: rd_data_1 <= 24'h7f007f;
		12'd1288: rd_data_1 <= 24'h7f007f;
		12'd1289: rd_data_1 <= 24'h7f007f;
		12'd1290: rd_data_1 <= 24'h7f007f;
		12'd1291: rd_data_1 <= 24'h7f007f;
		12'd1292: rd_data_1 <= 24'h7e007f;
		12'd1293: rd_data_1 <= 24'h7f007f;
		12'd1294: rd_data_1 <= 24'h7f007f;
		12'd1295: rd_data_1 <= 24'h80007d;
		12'd1296: rd_data_1 <= 24'h84007c;
		12'd1297: rd_data_1 <= 24'h83017c;
		12'd1298: rd_data_1 <= 24'h82017c;
		12'd1299: rd_data_1 <= 24'h81017a;
		12'd1300: rd_data_1 <= 24'h85057f;
		12'd1301: rd_data_1 <= 24'h81037b;
		12'd1302: rd_data_1 <= 24'h7d0077;
		12'd1303: rd_data_1 <= 24'h7f007a;
		12'd1304: rd_data_1 <= 24'h7e0079;
		12'd1305: rd_data_1 <= 24'h810081;
		12'd1306: rd_data_1 <= 24'h7e0081;
		12'd1307: rd_data_1 <= 24'h7e0184;
		12'd1308: rd_data_1 <= 24'h7e0086;
		12'd1309: rd_data_1 <= 24'h7e0084;
		12'd1310: rd_data_1 <= 24'h7e0082;
		12'd1311: rd_data_1 <= 24'h7c007d;
		12'd1312: rd_data_1 <= 24'h7c007f;
		12'd1313: rd_data_1 <= 24'h820385;
		12'd1314: rd_data_1 <= 24'h810483;
		12'd1315: rd_data_1 <= 24'h7e017e;
		12'd1316: rd_data_1 <= 24'h7f0181;
		12'd1317: rd_data_1 <= 24'h7d007e;
		12'd1318: rd_data_1 <= 24'h7d007e;
		12'd1319: rd_data_1 <= 24'h7d007d;
		12'd1320: rd_data_1 <= 24'h7d007c;
		12'd1321: rd_data_1 <= 24'h7e007c;
		12'd1322: rd_data_1 <= 24'h7e007d;
		12'd1323: rd_data_1 <= 24'h7e007e;
		12'd1324: rd_data_1 <= 24'h7e007e;
		12'd1325: rd_data_1 <= 24'h7e007e;
		12'd1326: rd_data_1 <= 24'h7e007e;
		12'd1327: rd_data_1 <= 24'h7e007e;
		12'd1328: rd_data_1 <= 24'h7e007e;
		12'd1329: rd_data_1 <= 24'h7f007f;
		12'd1330: rd_data_1 <= 24'h7f007f;
		12'd1331: rd_data_1 <= 24'h7f007f;
		12'd1332: rd_data_1 <= 24'h7f007f;
		12'd1333: rd_data_1 <= 24'h7f007f;
		12'd1334: rd_data_1 <= 24'h7f007f;
		12'd1335: rd_data_1 <= 24'h7f007f;
		12'd1336: rd_data_1 <= 24'h7f007f;
		12'd1337: rd_data_1 <= 24'h7f007f;
		12'd1338: rd_data_1 <= 24'h7f007f;
		12'd1339: rd_data_1 <= 24'h7f007f;
		12'd1340: rd_data_1 <= 24'h7f007f;
		12'd1341: rd_data_1 <= 24'h7f007f;
		12'd1342: rd_data_1 <= 24'h7f007f;
		12'd1343: rd_data_1 <= 24'h7f007f;
		12'd1344: rd_data_1 <= 24'h7f007f;
		12'd1345: rd_data_1 <= 24'h7f007f;
		12'd1346: rd_data_1 <= 24'h7f007f;
		12'd1347: rd_data_1 <= 24'h7f007f;
		12'd1348: rd_data_1 <= 24'h7f007f;
		12'd1349: rd_data_1 <= 24'h7f007f;
		12'd1350: rd_data_1 <= 24'h7f007f;
		12'd1351: rd_data_1 <= 24'h7f007f;
		12'd1352: rd_data_1 <= 24'h7f007f;
		12'd1353: rd_data_1 <= 24'h7f007f;
		12'd1354: rd_data_1 <= 24'h7f007f;
		12'd1355: rd_data_1 <= 24'h7f007f;
		12'd1356: rd_data_1 <= 24'h7f007f;
		12'd1357: rd_data_1 <= 24'h7f007f;
		12'd1358: rd_data_1 <= 24'h7f007d;
		12'd1359: rd_data_1 <= 24'h81007d;
		12'd1360: rd_data_1 <= 24'h82017c;
		12'd1361: rd_data_1 <= 24'h82017c;
		12'd1362: rd_data_1 <= 24'h82017c;
		12'd1363: rd_data_1 <= 24'h83007d;
		12'd1364: rd_data_1 <= 24'h84007e;
		12'd1365: rd_data_1 <= 24'h850080;
		12'd1366: rd_data_1 <= 24'h860081;
		12'd1367: rd_data_1 <= 24'h850081;
		12'd1368: rd_data_1 <= 24'h800082;
		12'd1369: rd_data_1 <= 24'h7b0181;
		12'd1370: rd_data_1 <= 24'h7e0080;
		12'd1371: rd_data_1 <= 24'h81007d;
		12'd1372: rd_data_1 <= 24'h81007c;
		12'd1373: rd_data_1 <= 24'h80007c;
		12'd1374: rd_data_1 <= 24'h7f007f;
		12'd1375: rd_data_1 <= 24'h7d007f;
		12'd1376: rd_data_1 <= 24'h7c017c;
		12'd1377: rd_data_1 <= 24'h7c0377;
		12'd1378: rd_data_1 <= 24'h7c0377;
		12'd1379: rd_data_1 <= 24'h7d0278;
		12'd1380: rd_data_1 <= 24'h7e0279;
		12'd1381: rd_data_1 <= 24'h7e017c;
		12'd1382: rd_data_1 <= 24'h7e017e;
		12'd1383: rd_data_1 <= 24'h7e007f;
		12'd1384: rd_data_1 <= 24'h7e007f;
		12'd1385: rd_data_1 <= 24'h7f007f;
		12'd1386: rd_data_1 <= 24'h7f007f;
		12'd1387: rd_data_1 <= 24'h7f007f;
		12'd1388: rd_data_1 <= 24'h7f007f;
		12'd1389: rd_data_1 <= 24'h7f007f;
		12'd1390: rd_data_1 <= 24'h7f007f;
		12'd1391: rd_data_1 <= 24'h7f007f;
		12'd1392: rd_data_1 <= 24'h7f007f;
		12'd1393: rd_data_1 <= 24'h7f007f;
		12'd1394: rd_data_1 <= 24'h7f007f;
		12'd1395: rd_data_1 <= 24'h7f007f;
		12'd1396: rd_data_1 <= 24'h7f007f;
		12'd1397: rd_data_1 <= 24'h7f007f;
		12'd1398: rd_data_1 <= 24'h7f007f;
		12'd1399: rd_data_1 <= 24'h7f007f;
		12'd1400: rd_data_1 <= 24'h7f007f;
		12'd1401: rd_data_1 <= 24'h7f007f;
		12'd1402: rd_data_1 <= 24'h7f007f;
		12'd1403: rd_data_1 <= 24'h7f007f;
		12'd1404: rd_data_1 <= 24'h7f007f;
		12'd1405: rd_data_1 <= 24'h7f007f;
		12'd1406: rd_data_1 <= 24'h7f007f;
		12'd1407: rd_data_1 <= 24'h7f007f;
		12'd1408: rd_data_1 <= 24'h7f007f;
		12'd1409: rd_data_1 <= 24'h7f007f;
		12'd1410: rd_data_1 <= 24'h7f007f;
		12'd1411: rd_data_1 <= 24'h7f007f;
		12'd1412: rd_data_1 <= 24'h7f007f;
		12'd1413: rd_data_1 <= 24'h7f007f;
		12'd1414: rd_data_1 <= 24'h7f007f;
		12'd1415: rd_data_1 <= 24'h7f007f;
		12'd1416: rd_data_1 <= 24'h7f007f;
		12'd1417: rd_data_1 <= 24'h7f007f;
		12'd1418: rd_data_1 <= 24'h7f007f;
		12'd1419: rd_data_1 <= 24'h7f007f;
		12'd1420: rd_data_1 <= 24'h7f007f;
		12'd1421: rd_data_1 <= 24'h7f007f;
		12'd1422: rd_data_1 <= 24'h7f007d;
		12'd1423: rd_data_1 <= 24'h7f007d;
		12'd1424: rd_data_1 <= 24'h810080;
		12'd1425: rd_data_1 <= 24'h820081;
		12'd1426: rd_data_1 <= 24'h820081;
		12'd1427: rd_data_1 <= 24'h830081;
		12'd1428: rd_data_1 <= 24'h840081;
		12'd1429: rd_data_1 <= 24'h840082;
		12'd1430: rd_data_1 <= 24'h840082;
		12'd1431: rd_data_1 <= 24'h830082;
		12'd1432: rd_data_1 <= 24'h7d0182;
		12'd1433: rd_data_1 <= 24'h7a0280;
		12'd1434: rd_data_1 <= 24'h7d017e;
		12'd1435: rd_data_1 <= 24'h80007d;
		12'd1436: rd_data_1 <= 24'h80007d;
		12'd1437: rd_data_1 <= 24'h7e007c;
		12'd1438: rd_data_1 <= 24'h7b007d;
		12'd1439: rd_data_1 <= 24'h7a007d;
		12'd1440: rd_data_1 <= 24'h7c027a;
		12'd1441: rd_data_1 <= 24'h800276;
		12'd1442: rd_data_1 <= 24'h800275;
		12'd1443: rd_data_1 <= 24'h800276;
		12'd1444: rd_data_1 <= 24'h7f0079;
		12'd1445: rd_data_1 <= 24'h7f007c;
		12'd1446: rd_data_1 <= 24'h7e017d;
		12'd1447: rd_data_1 <= 24'h7e017e;
		12'd1448: rd_data_1 <= 24'h7e007f;
		12'd1449: rd_data_1 <= 24'h7f007f;
		12'd1450: rd_data_1 <= 24'h7f007f;
		12'd1451: rd_data_1 <= 24'h7f007f;
		12'd1452: rd_data_1 <= 24'h7f007f;
		12'd1453: rd_data_1 <= 24'h7f007f;
		12'd1454: rd_data_1 <= 24'h7f007f;
		12'd1455: rd_data_1 <= 24'h7f007f;
		12'd1456: rd_data_1 <= 24'h7f007f;
		12'd1457: rd_data_1 <= 24'h7f007f;
		12'd1458: rd_data_1 <= 24'h7f007f;
		12'd1459: rd_data_1 <= 24'h7f007f;
		12'd1460: rd_data_1 <= 24'h7f007f;
		12'd1461: rd_data_1 <= 24'h7f007f;
		12'd1462: rd_data_1 <= 24'h7f007f;
		12'd1463: rd_data_1 <= 24'h7f007f;
		12'd1464: rd_data_1 <= 24'h7f007f;
		12'd1465: rd_data_1 <= 24'h7f007f;
		12'd1466: rd_data_1 <= 24'h7f007f;
		12'd1467: rd_data_1 <= 24'h7f007f;
		12'd1468: rd_data_1 <= 24'h7f007f;
		12'd1469: rd_data_1 <= 24'h7f007f;
		12'd1470: rd_data_1 <= 24'h7f007f;
		12'd1471: rd_data_1 <= 24'h7f007f;
		12'd1472: rd_data_1 <= 24'h7f007f;
		12'd1473: rd_data_1 <= 24'h7f007f;
		12'd1474: rd_data_1 <= 24'h7f007f;
		12'd1475: rd_data_1 <= 24'h7f007f;
		12'd1476: rd_data_1 <= 24'h7f007f;
		12'd1477: rd_data_1 <= 24'h7f007f;
		12'd1478: rd_data_1 <= 24'h7f007f;
		12'd1479: rd_data_1 <= 24'h7f007f;
		12'd1480: rd_data_1 <= 24'h7f007f;
		12'd1481: rd_data_1 <= 24'h7f007f;
		12'd1482: rd_data_1 <= 24'h7f007f;
		12'd1483: rd_data_1 <= 24'h7f007f;
		12'd1484: rd_data_1 <= 24'h7f007f;
		12'd1485: rd_data_1 <= 24'h7f007f;
		12'd1486: rd_data_1 <= 24'h81007f;
		12'd1487: rd_data_1 <= 24'h810080;
		12'd1488: rd_data_1 <= 24'h820085;
		12'd1489: rd_data_1 <= 24'h820088;
		12'd1490: rd_data_1 <= 24'h820087;
		12'd1491: rd_data_1 <= 24'h810085;
		12'd1492: rd_data_1 <= 24'h800182;
		12'd1493: rd_data_1 <= 24'h7e0182;
		12'd1494: rd_data_1 <= 24'h7d0281;
		12'd1495: rd_data_1 <= 24'h7d0280;
		12'd1496: rd_data_1 <= 24'h7c027e;
		12'd1497: rd_data_1 <= 24'h7d017d;
		12'd1498: rd_data_1 <= 24'h7e007f;
		12'd1499: rd_data_1 <= 24'h7e0082;
		12'd1500: rd_data_1 <= 24'h7c0083;
		12'd1501: rd_data_1 <= 24'h7a0081;
		12'd1502: rd_data_1 <= 24'h77027e;
		12'd1503: rd_data_1 <= 24'h77037b;
		12'd1504: rd_data_1 <= 24'h7e0179;
		12'd1505: rd_data_1 <= 24'h880079;
		12'd1506: rd_data_1 <= 24'h89007a;
		12'd1507: rd_data_1 <= 24'h86007a;
		12'd1508: rd_data_1 <= 24'h83007b;
		12'd1509: rd_data_1 <= 24'h80007c;
		12'd1510: rd_data_1 <= 24'h7e007d;
		12'd1511: rd_data_1 <= 24'h7e017d;
		12'd1512: rd_data_1 <= 24'h7e017e;
		12'd1513: rd_data_1 <= 24'h7f007f;
		12'd1514: rd_data_1 <= 24'h7f007f;
		12'd1515: rd_data_1 <= 24'h7f007f;
		12'd1516: rd_data_1 <= 24'h7f007f;
		12'd1517: rd_data_1 <= 24'h7f007f;
		12'd1518: rd_data_1 <= 24'h7f007f;
		12'd1519: rd_data_1 <= 24'h7f007f;
		12'd1520: rd_data_1 <= 24'h7f007f;
		12'd1521: rd_data_1 <= 24'h7f007f;
		12'd1522: rd_data_1 <= 24'h7f007f;
		12'd1523: rd_data_1 <= 24'h7f007f;
		12'd1524: rd_data_1 <= 24'h7f007f;
		12'd1525: rd_data_1 <= 24'h7f007f;
		12'd1526: rd_data_1 <= 24'h7f007f;
		12'd1527: rd_data_1 <= 24'h7f007f;
		12'd1528: rd_data_1 <= 24'h7f007f;
		12'd1529: rd_data_1 <= 24'h7f007f;
		12'd1530: rd_data_1 <= 24'h7f007f;
		12'd1531: rd_data_1 <= 24'h7f007f;
		12'd1532: rd_data_1 <= 24'h7f007f;
		12'd1533: rd_data_1 <= 24'h7f007f;
		12'd1534: rd_data_1 <= 24'h7f007f;
		12'd1535: rd_data_1 <= 24'h7f007f;
		12'd1536: rd_data_1 <= 24'h7f007f;
		12'd1537: rd_data_1 <= 24'h7f007f;
		12'd1538: rd_data_1 <= 24'h7f007f;
		12'd1539: rd_data_1 <= 24'h7f007f;
		12'd1540: rd_data_1 <= 24'h7f007f;
		12'd1541: rd_data_1 <= 24'h7f007f;
		12'd1542: rd_data_1 <= 24'h7f007f;
		12'd1543: rd_data_1 <= 24'h7f007f;
		12'd1544: rd_data_1 <= 24'h7f007f;
		12'd1545: rd_data_1 <= 24'h7f007f;
		12'd1546: rd_data_1 <= 24'h7f007f;
		12'd1547: rd_data_1 <= 24'h7f007f;
		12'd1548: rd_data_1 <= 24'h7f007f;
		12'd1549: rd_data_1 <= 24'h7f007f;
		12'd1550: rd_data_1 <= 24'h81007f;
		12'd1551: rd_data_1 <= 24'h810080;
		12'd1552: rd_data_1 <= 24'h820085;
		12'd1553: rd_data_1 <= 24'h820088;
		12'd1554: rd_data_1 <= 24'h810087;
		12'd1555: rd_data_1 <= 24'h800185;
		12'd1556: rd_data_1 <= 24'h7e0283;
		12'd1557: rd_data_1 <= 24'h7c0381;
		12'd1558: rd_data_1 <= 24'h7c0380;
		12'd1559: rd_data_1 <= 24'h7c047f;
		12'd1560: rd_data_1 <= 24'h7d027d;
		12'd1561: rd_data_1 <= 24'h7f007d;
		12'd1562: rd_data_1 <= 24'h7e007f;
		12'd1563: rd_data_1 <= 24'h7e0082;
		12'd1564: rd_data_1 <= 24'h7d0083;
		12'd1565: rd_data_1 <= 24'h790081;
		12'd1566: rd_data_1 <= 24'h76027e;
		12'd1567: rd_data_1 <= 24'h78027c;
		12'd1568: rd_data_1 <= 24'h81007c;
		12'd1569: rd_data_1 <= 24'h88007d;
		12'd1570: rd_data_1 <= 24'h88007d;
		12'd1571: rd_data_1 <= 24'h87007d;
		12'd1572: rd_data_1 <= 24'h85007d;
		12'd1573: rd_data_1 <= 24'h81007d;
		12'd1574: rd_data_1 <= 24'h7e007d;
		12'd1575: rd_data_1 <= 24'h7e017d;
		12'd1576: rd_data_1 <= 24'h7e017e;
		12'd1577: rd_data_1 <= 24'h7f007f;
		12'd1578: rd_data_1 <= 24'h7f007f;
		12'd1579: rd_data_1 <= 24'h7f007f;
		12'd1580: rd_data_1 <= 24'h7f007f;
		12'd1581: rd_data_1 <= 24'h7f007f;
		12'd1582: rd_data_1 <= 24'h7f007f;
		12'd1583: rd_data_1 <= 24'h7f007f;
		12'd1584: rd_data_1 <= 24'h7f007f;
		12'd1585: rd_data_1 <= 24'h7f007f;
		12'd1586: rd_data_1 <= 24'h7f007f;
		12'd1587: rd_data_1 <= 24'h7f007f;
		12'd1588: rd_data_1 <= 24'h7f007f;
		12'd1589: rd_data_1 <= 24'h7f007f;
		12'd1590: rd_data_1 <= 24'h7f007f;
		12'd1591: rd_data_1 <= 24'h7f007f;
		12'd1592: rd_data_1 <= 24'h7f007f;
		12'd1593: rd_data_1 <= 24'h7f007f;
		12'd1594: rd_data_1 <= 24'h7f007f;
		12'd1595: rd_data_1 <= 24'h7f007f;
		12'd1596: rd_data_1 <= 24'h7f007f;
		12'd1597: rd_data_1 <= 24'h7f007f;
		12'd1598: rd_data_1 <= 24'h7f007f;
		12'd1599: rd_data_1 <= 24'h7f007f;
		12'd1600: rd_data_1 <= 24'h7f007f;
		12'd1601: rd_data_1 <= 24'h7f007f;
		12'd1602: rd_data_1 <= 24'h7f007f;
		12'd1603: rd_data_1 <= 24'h7f007f;
		12'd1604: rd_data_1 <= 24'h7f007f;
		12'd1605: rd_data_1 <= 24'h7f007f;
		12'd1606: rd_data_1 <= 24'h7f007f;
		12'd1607: rd_data_1 <= 24'h7f007f;
		12'd1608: rd_data_1 <= 24'h7f007f;
		12'd1609: rd_data_1 <= 24'h7f007f;
		12'd1610: rd_data_1 <= 24'h7f007f;
		12'd1611: rd_data_1 <= 24'h7f007f;
		12'd1612: rd_data_1 <= 24'h7f007f;
		12'd1613: rd_data_1 <= 24'h7f007f;
		12'd1614: rd_data_1 <= 24'h7f007f;
		12'd1615: rd_data_1 <= 24'h7f007f;
		12'd1616: rd_data_1 <= 24'h810081;
		12'd1617: rd_data_1 <= 24'h810082;
		12'd1618: rd_data_1 <= 24'h810082;
		12'd1619: rd_data_1 <= 24'h810082;
		12'd1620: rd_data_1 <= 24'h800181;
		12'd1621: rd_data_1 <= 24'h7f0280;
		12'd1622: rd_data_1 <= 24'h7f0280;
		12'd1623: rd_data_1 <= 24'h7f0280;
		12'd1624: rd_data_1 <= 24'h800180;
		12'd1625: rd_data_1 <= 24'h810180;
		12'd1626: rd_data_1 <= 24'h810180;
		12'd1627: rd_data_1 <= 24'h810081;
		12'd1628: rd_data_1 <= 24'h7f0082;
		12'd1629: rd_data_1 <= 24'h7e0080;
		12'd1630: rd_data_1 <= 24'h7d017f;
		12'd1631: rd_data_1 <= 24'h7d017f;
		12'd1632: rd_data_1 <= 24'h7f007f;
		12'd1633: rd_data_1 <= 24'h82007f;
		12'd1634: rd_data_1 <= 24'h83007f;
		12'd1635: rd_data_1 <= 24'h82007f;
		12'd1636: rd_data_1 <= 24'h81007f;
		12'd1637: rd_data_1 <= 24'h80007f;
		12'd1638: rd_data_1 <= 24'h7f007f;
		12'd1639: rd_data_1 <= 24'h7f007f;
		12'd1640: rd_data_1 <= 24'h7f007f;
		12'd1641: rd_data_1 <= 24'h7f007f;
		12'd1642: rd_data_1 <= 24'h7f007f;
		12'd1643: rd_data_1 <= 24'h7f007f;
		12'd1644: rd_data_1 <= 24'h7f007f;
		12'd1645: rd_data_1 <= 24'h7f007f;
		12'd1646: rd_data_1 <= 24'h7f007f;
		12'd1647: rd_data_1 <= 24'h7f007f;
		12'd1648: rd_data_1 <= 24'h7f007f;
		12'd1649: rd_data_1 <= 24'h7f007f;
		12'd1650: rd_data_1 <= 24'h7f007f;
		12'd1651: rd_data_1 <= 24'h7f007f;
		12'd1652: rd_data_1 <= 24'h7f007f;
		12'd1653: rd_data_1 <= 24'h7f007f;
		12'd1654: rd_data_1 <= 24'h7f007f;
		12'd1655: rd_data_1 <= 24'h7f007f;
		12'd1656: rd_data_1 <= 24'h7f007f;
		12'd1657: rd_data_1 <= 24'h7f007f;
		12'd1658: rd_data_1 <= 24'h7f007f;
		12'd1659: rd_data_1 <= 24'h7f007f;
		12'd1660: rd_data_1 <= 24'h7f007f;
		12'd1661: rd_data_1 <= 24'h7f007f;
		12'd1662: rd_data_1 <= 24'h7f007f;
		12'd1663: rd_data_1 <= 24'h7f007f;
		12'd1664: rd_data_1 <= 24'h7f007f;
		12'd1665: rd_data_1 <= 24'h7f007f;
		12'd1666: rd_data_1 <= 24'h7f007f;
		12'd1667: rd_data_1 <= 24'h7f007f;
		12'd1668: rd_data_1 <= 24'h7f007f;
		12'd1669: rd_data_1 <= 24'h7f007f;
		12'd1670: rd_data_1 <= 24'h7f007f;
		12'd1671: rd_data_1 <= 24'h7f007f;
		12'd1672: rd_data_1 <= 24'h7f007f;
		12'd1673: rd_data_1 <= 24'h7f007f;
		12'd1674: rd_data_1 <= 24'h7f007f;
		12'd1675: rd_data_1 <= 24'h7f007f;
		12'd1676: rd_data_1 <= 24'h7f007f;
		12'd1677: rd_data_1 <= 24'h7f007f;
		12'd1678: rd_data_1 <= 24'h7f007f;
		12'd1679: rd_data_1 <= 24'h7f007f;
		12'd1680: rd_data_1 <= 24'h810180;
		12'd1681: rd_data_1 <= 24'h810180;
		12'd1682: rd_data_1 <= 24'h810180;
		12'd1683: rd_data_1 <= 24'h810180;
		12'd1684: rd_data_1 <= 24'h810180;
		12'd1685: rd_data_1 <= 24'h810180;
		12'd1686: rd_data_1 <= 24'h810180;
		12'd1687: rd_data_1 <= 24'h810180;
		12'd1688: rd_data_1 <= 24'h810180;
		12'd1689: rd_data_1 <= 24'h810180;
		12'd1690: rd_data_1 <= 24'h810180;
		12'd1691: rd_data_1 <= 24'h810180;
		12'd1692: rd_data_1 <= 24'h80007f;
		12'd1693: rd_data_1 <= 24'h7f007f;
		12'd1694: rd_data_1 <= 24'h7f007f;
		12'd1695: rd_data_1 <= 24'h7f007f;
		12'd1696: rd_data_1 <= 24'h7f007f;
		12'd1697: rd_data_1 <= 24'h7f007f;
		12'd1698: rd_data_1 <= 24'h7f007f;
		12'd1699: rd_data_1 <= 24'h7f007f;
		12'd1700: rd_data_1 <= 24'h7f007f;
		12'd1701: rd_data_1 <= 24'h7f007f;
		12'd1702: rd_data_1 <= 24'h7f007f;
		12'd1703: rd_data_1 <= 24'h7f007f;
		12'd1704: rd_data_1 <= 24'h7f007f;
		12'd1705: rd_data_1 <= 24'h7f007f;
		12'd1706: rd_data_1 <= 24'h7f007f;
		12'd1707: rd_data_1 <= 24'h7f007f;
		12'd1708: rd_data_1 <= 24'h7f007f;
		12'd1709: rd_data_1 <= 24'h7f007f;
		12'd1710: rd_data_1 <= 24'h7f007f;
		12'd1711: rd_data_1 <= 24'h7f007f;
		12'd1712: rd_data_1 <= 24'h7f007f;
		12'd1713: rd_data_1 <= 24'h7f007f;
		12'd1714: rd_data_1 <= 24'h7f007f;
		12'd1715: rd_data_1 <= 24'h7f007f;
		12'd1716: rd_data_1 <= 24'h7f007f;
		12'd1717: rd_data_1 <= 24'h7f007f;
		12'd1718: rd_data_1 <= 24'h7f007f;
		12'd1719: rd_data_1 <= 24'h7f007f;
		12'd1720: rd_data_1 <= 24'h7f007f;
		12'd1721: rd_data_1 <= 24'h7f007f;
		12'd1722: rd_data_1 <= 24'h7f007f;
		12'd1723: rd_data_1 <= 24'h7f007f;
		12'd1724: rd_data_1 <= 24'h7f007f;
		12'd1725: rd_data_1 <= 24'h7f007f;
		12'd1726: rd_data_1 <= 24'h7f007f;
		12'd1727: rd_data_1 <= 24'h7f007f;
		12'd1728: rd_data_1 <= 24'h7f007f;
		12'd1729: rd_data_1 <= 24'h7f007f;
		12'd1730: rd_data_1 <= 24'h7f007f;
		12'd1731: rd_data_1 <= 24'h7f007f;
		12'd1732: rd_data_1 <= 24'h7f007f;
		12'd1733: rd_data_1 <= 24'h7f007f;
		12'd1734: rd_data_1 <= 24'h7f007f;
		12'd1735: rd_data_1 <= 24'h7f007f;
		12'd1736: rd_data_1 <= 24'h7f007f;
		12'd1737: rd_data_1 <= 24'h7f007f;
		12'd1738: rd_data_1 <= 24'h7f007f;
		12'd1739: rd_data_1 <= 24'h7f007f;
		12'd1740: rd_data_1 <= 24'h7f007f;
		12'd1741: rd_data_1 <= 24'h7f007f;
		12'd1742: rd_data_1 <= 24'h7f007f;
		12'd1743: rd_data_1 <= 24'h7f007f;
		12'd1744: rd_data_1 <= 24'h810180;
		12'd1745: rd_data_1 <= 24'h810180;
		12'd1746: rd_data_1 <= 24'h810180;
		12'd1747: rd_data_1 <= 24'h810180;
		12'd1748: rd_data_1 <= 24'h810180;
		12'd1749: rd_data_1 <= 24'h810180;
		12'd1750: rd_data_1 <= 24'h810180;
		12'd1751: rd_data_1 <= 24'h810180;
		12'd1752: rd_data_1 <= 24'h810180;
		12'd1753: rd_data_1 <= 24'h810180;
		12'd1754: rd_data_1 <= 24'h810180;
		12'd1755: rd_data_1 <= 24'h810180;
		12'd1756: rd_data_1 <= 24'h80007f;
		12'd1757: rd_data_1 <= 24'h7f007f;
		12'd1758: rd_data_1 <= 24'h7f007f;
		12'd1759: rd_data_1 <= 24'h7f007f;
		12'd1760: rd_data_1 <= 24'h7f007f;
		12'd1761: rd_data_1 <= 24'h7f007f;
		12'd1762: rd_data_1 <= 24'h7f007f;
		12'd1763: rd_data_1 <= 24'h7f007f;
		12'd1764: rd_data_1 <= 24'h7f007f;
		12'd1765: rd_data_1 <= 24'h7f007f;
		12'd1766: rd_data_1 <= 24'h7f007f;
		12'd1767: rd_data_1 <= 24'h7f007f;
		12'd1768: rd_data_1 <= 24'h7f007f;
		12'd1769: rd_data_1 <= 24'h7f007f;
		12'd1770: rd_data_1 <= 24'h7f007f;
		12'd1771: rd_data_1 <= 24'h7f007f;
		12'd1772: rd_data_1 <= 24'h7f007f;
		12'd1773: rd_data_1 <= 24'h7f007f;
		12'd1774: rd_data_1 <= 24'h7f007f;
		12'd1775: rd_data_1 <= 24'h7f007f;
		12'd1776: rd_data_1 <= 24'h7f007f;
		12'd1777: rd_data_1 <= 24'h7f007f;
		12'd1778: rd_data_1 <= 24'h7f007f;
		12'd1779: rd_data_1 <= 24'h7f007f;
		12'd1780: rd_data_1 <= 24'h7f007f;
		12'd1781: rd_data_1 <= 24'h7f007f;
		12'd1782: rd_data_1 <= 24'h7f007f;
		12'd1783: rd_data_1 <= 24'h7f007f;
		12'd1784: rd_data_1 <= 24'h7f007f;
		12'd1785: rd_data_1 <= 24'h7f007f;
		12'd1786: rd_data_1 <= 24'h7f007f;
		12'd1787: rd_data_1 <= 24'h7f007f;
		12'd1788: rd_data_1 <= 24'h7f007f;
		12'd1789: rd_data_1 <= 24'h7f007f;
		12'd1790: rd_data_1 <= 24'h7f007f;
		12'd1791: rd_data_1 <= 24'h7f007f;
		12'd1792: rd_data_1 <= 24'h7f007f;
		12'd1793: rd_data_1 <= 24'h7f007f;
		12'd1794: rd_data_1 <= 24'h7f007f;
		12'd1795: rd_data_1 <= 24'h7f007f;
		12'd1796: rd_data_1 <= 24'h7f007f;
		12'd1797: rd_data_1 <= 24'h7f007f;
		12'd1798: rd_data_1 <= 24'h7f007f;
		12'd1799: rd_data_1 <= 24'h7f007f;
		12'd1800: rd_data_1 <= 24'h7f007f;
		12'd1801: rd_data_1 <= 24'h7f007f;
		12'd1802: rd_data_1 <= 24'h7f007f;
		12'd1803: rd_data_1 <= 24'h7f007f;
		12'd1804: rd_data_1 <= 24'h7f007f;
		12'd1805: rd_data_1 <= 24'h7f007f;
		12'd1806: rd_data_1 <= 24'h7f007f;
		12'd1807: rd_data_1 <= 24'h7f007f;
		12'd1808: rd_data_1 <= 24'h810180;
		12'd1809: rd_data_1 <= 24'h810180;
		12'd1810: rd_data_1 <= 24'h810180;
		12'd1811: rd_data_1 <= 24'h810180;
		12'd1812: rd_data_1 <= 24'h810180;
		12'd1813: rd_data_1 <= 24'h810180;
		12'd1814: rd_data_1 <= 24'h810180;
		12'd1815: rd_data_1 <= 24'h810180;
		12'd1816: rd_data_1 <= 24'h810180;
		12'd1817: rd_data_1 <= 24'h810180;
		12'd1818: rd_data_1 <= 24'h810180;
		12'd1819: rd_data_1 <= 24'h810180;
		12'd1820: rd_data_1 <= 24'h80007f;
		12'd1821: rd_data_1 <= 24'h7f007f;
		12'd1822: rd_data_1 <= 24'h7f007f;
		12'd1823: rd_data_1 <= 24'h7f007f;
		12'd1824: rd_data_1 <= 24'h7f007f;
		12'd1825: rd_data_1 <= 24'h7f007f;
		12'd1826: rd_data_1 <= 24'h7f007f;
		12'd1827: rd_data_1 <= 24'h7f007f;
		12'd1828: rd_data_1 <= 24'h7f007f;
		12'd1829: rd_data_1 <= 24'h7f007f;
		12'd1830: rd_data_1 <= 24'h7f007f;
		12'd1831: rd_data_1 <= 24'h7f007f;
		12'd1832: rd_data_1 <= 24'h7f007f;
		12'd1833: rd_data_1 <= 24'h7f007f;
		12'd1834: rd_data_1 <= 24'h7f007f;
		12'd1835: rd_data_1 <= 24'h7f007f;
		12'd1836: rd_data_1 <= 24'h7f007f;
		12'd1837: rd_data_1 <= 24'h7f007f;
		12'd1838: rd_data_1 <= 24'h7f007f;
		12'd1839: rd_data_1 <= 24'h7f007f;
		12'd1840: rd_data_1 <= 24'h7f007f;
		12'd1841: rd_data_1 <= 24'h7f007f;
		12'd1842: rd_data_1 <= 24'h7f007f;
		12'd1843: rd_data_1 <= 24'h7f007f;
		12'd1844: rd_data_1 <= 24'h7f007f;
		12'd1845: rd_data_1 <= 24'h7f007f;
		12'd1846: rd_data_1 <= 24'h7f007f;
		12'd1847: rd_data_1 <= 24'h7f007f;
		12'd1848: rd_data_1 <= 24'h7f007f;
		12'd1849: rd_data_1 <= 24'h7f007f;
		12'd1850: rd_data_1 <= 24'h7f007f;
		12'd1851: rd_data_1 <= 24'h7f007f;
		12'd1852: rd_data_1 <= 24'h7f007f;
		12'd1853: rd_data_1 <= 24'h7f007f;
		12'd1854: rd_data_1 <= 24'h7f007f;
		12'd1855: rd_data_1 <= 24'h7f007f;
		12'd1856: rd_data_1 <= 24'h7f007f;
		12'd1857: rd_data_1 <= 24'h7f007f;
		12'd1858: rd_data_1 <= 24'h7f007f;
		12'd1859: rd_data_1 <= 24'h7f007f;
		12'd1860: rd_data_1 <= 24'h7f007f;
		12'd1861: rd_data_1 <= 24'h7f007f;
		12'd1862: rd_data_1 <= 24'h7f007f;
		12'd1863: rd_data_1 <= 24'h7f007f;
		12'd1864: rd_data_1 <= 24'h7f007f;
		12'd1865: rd_data_1 <= 24'h7f007f;
		12'd1866: rd_data_1 <= 24'h7f007f;
		12'd1867: rd_data_1 <= 24'h7f007f;
		12'd1868: rd_data_1 <= 24'h7f007f;
		12'd1869: rd_data_1 <= 24'h7f007f;
		12'd1870: rd_data_1 <= 24'h7f007f;
		12'd1871: rd_data_1 <= 24'h7f007f;
		12'd1872: rd_data_1 <= 24'h810180;
		12'd1873: rd_data_1 <= 24'h810180;
		12'd1874: rd_data_1 <= 24'h810180;
		12'd1875: rd_data_1 <= 24'h810180;
		12'd1876: rd_data_1 <= 24'h810180;
		12'd1877: rd_data_1 <= 24'h810180;
		12'd1878: rd_data_1 <= 24'h810180;
		12'd1879: rd_data_1 <= 24'h810180;
		12'd1880: rd_data_1 <= 24'h810180;
		12'd1881: rd_data_1 <= 24'h810180;
		12'd1882: rd_data_1 <= 24'h810180;
		12'd1883: rd_data_1 <= 24'h810180;
		12'd1884: rd_data_1 <= 24'h810180;
		12'd1885: rd_data_1 <= 24'h810180;
		12'd1886: rd_data_1 <= 24'h810180;
		12'd1887: rd_data_1 <= 24'h810180;
		12'd1888: rd_data_1 <= 24'h810180;
		12'd1889: rd_data_1 <= 24'h810180;
		12'd1890: rd_data_1 <= 24'h810180;
		12'd1891: rd_data_1 <= 24'h810180;
		12'd1892: rd_data_1 <= 24'h810180;
		12'd1893: rd_data_1 <= 24'h810180;
		12'd1894: rd_data_1 <= 24'h810180;
		12'd1895: rd_data_1 <= 24'h810180;
		12'd1896: rd_data_1 <= 24'h810180;
		12'd1897: rd_data_1 <= 24'h810180;
		12'd1898: rd_data_1 <= 24'h810180;
		12'd1899: rd_data_1 <= 24'h810180;
		12'd1900: rd_data_1 <= 24'h810180;
		12'd1901: rd_data_1 <= 24'h810180;
		12'd1902: rd_data_1 <= 24'h810180;
		12'd1903: rd_data_1 <= 24'h810180;
		12'd1904: rd_data_1 <= 24'h810180;
		12'd1905: rd_data_1 <= 24'h7f007f;
		12'd1906: rd_data_1 <= 24'h7f007f;
		12'd1907: rd_data_1 <= 24'h7f007f;
		12'd1908: rd_data_1 <= 24'h7f007f;
		12'd1909: rd_data_1 <= 24'h7f007f;
		12'd1910: rd_data_1 <= 24'h7f007f;
		12'd1911: rd_data_1 <= 24'h7f007f;
		12'd1912: rd_data_1 <= 24'h7f007f;
		12'd1913: rd_data_1 <= 24'h7f007f;
		12'd1914: rd_data_1 <= 24'h7f007f;
		12'd1915: rd_data_1 <= 24'h7f007f;
		12'd1916: rd_data_1 <= 24'h7f007f;
		12'd1917: rd_data_1 <= 24'h7f007f;
		12'd1918: rd_data_1 <= 24'h7f007f;
		12'd1919: rd_data_1 <= 24'h7f007f;
		12'd1920: rd_data_1 <= 24'h7f007f;
		12'd1921: rd_data_1 <= 24'h7f007f;
		12'd1922: rd_data_1 <= 24'h7f007f;
		12'd1923: rd_data_1 <= 24'h7f007f;
		12'd1924: rd_data_1 <= 24'h7f007f;
		12'd1925: rd_data_1 <= 24'h7f007f;
		12'd1926: rd_data_1 <= 24'h7f007f;
		12'd1927: rd_data_1 <= 24'h7f007f;
		12'd1928: rd_data_1 <= 24'h7f007f;
		12'd1929: rd_data_1 <= 24'h7f007f;
		12'd1930: rd_data_1 <= 24'h7f007f;
		12'd1931: rd_data_1 <= 24'h7f007f;
		12'd1932: rd_data_1 <= 24'h7f007f;
		12'd1933: rd_data_1 <= 24'h7f007f;
		12'd1934: rd_data_1 <= 24'h7f007f;
		12'd1935: rd_data_1 <= 24'h7f007f;
		12'd1936: rd_data_1 <= 24'h810180;
		12'd1937: rd_data_1 <= 24'h810180;
		12'd1938: rd_data_1 <= 24'h810180;
		12'd1939: rd_data_1 <= 24'h810180;
		12'd1940: rd_data_1 <= 24'h810180;
		12'd1941: rd_data_1 <= 24'h810180;
		12'd1942: rd_data_1 <= 24'h810180;
		12'd1943: rd_data_1 <= 24'h810180;
		12'd1944: rd_data_1 <= 24'h810180;
		12'd1945: rd_data_1 <= 24'h810180;
		12'd1946: rd_data_1 <= 24'h810180;
		12'd1947: rd_data_1 <= 24'h810180;
		12'd1948: rd_data_1 <= 24'h810180;
		12'd1949: rd_data_1 <= 24'h810180;
		12'd1950: rd_data_1 <= 24'h810180;
		12'd1951: rd_data_1 <= 24'h810180;
		12'd1952: rd_data_1 <= 24'h810180;
		12'd1953: rd_data_1 <= 24'h810180;
		12'd1954: rd_data_1 <= 24'h810180;
		12'd1955: rd_data_1 <= 24'h810180;
		12'd1956: rd_data_1 <= 24'h810180;
		12'd1957: rd_data_1 <= 24'h810180;
		12'd1958: rd_data_1 <= 24'h810180;
		12'd1959: rd_data_1 <= 24'h810180;
		12'd1960: rd_data_1 <= 24'h810180;
		12'd1961: rd_data_1 <= 24'h810180;
		12'd1962: rd_data_1 <= 24'h810180;
		12'd1963: rd_data_1 <= 24'h810180;
		12'd1964: rd_data_1 <= 24'h810180;
		12'd1965: rd_data_1 <= 24'h810180;
		12'd1966: rd_data_1 <= 24'h810180;
		12'd1967: rd_data_1 <= 24'h810180;
		12'd1968: rd_data_1 <= 24'h810180;
		12'd1969: rd_data_1 <= 24'h7f007f;
		12'd1970: rd_data_1 <= 24'h7f007f;
		12'd1971: rd_data_1 <= 24'h7f007f;
		12'd1972: rd_data_1 <= 24'h7f007f;
		12'd1973: rd_data_1 <= 24'h7f007f;
		12'd1974: rd_data_1 <= 24'h7f007f;
		12'd1975: rd_data_1 <= 24'h7f007f;
		12'd1976: rd_data_1 <= 24'h7f007f;
		12'd1977: rd_data_1 <= 24'h7f007f;
		12'd1978: rd_data_1 <= 24'h7f007f;
		12'd1979: rd_data_1 <= 24'h7f007f;
		12'd1980: rd_data_1 <= 24'h7f007f;
		12'd1981: rd_data_1 <= 24'h7f007f;
		12'd1982: rd_data_1 <= 24'h7f007f;
		12'd1983: rd_data_1 <= 24'h7f007f;
		12'd1984: rd_data_1 <= 24'h7f007f;
		12'd1985: rd_data_1 <= 24'h7f007f;
		12'd1986: rd_data_1 <= 24'h7f007f;
		12'd1987: rd_data_1 <= 24'h7f007f;
		12'd1988: rd_data_1 <= 24'h7f007f;
		12'd1989: rd_data_1 <= 24'h7f007f;
		12'd1990: rd_data_1 <= 24'h7f007f;
		12'd1991: rd_data_1 <= 24'h7f007f;
		12'd1992: rd_data_1 <= 24'h7f007f;
		12'd1993: rd_data_1 <= 24'h7f007f;
		12'd1994: rd_data_1 <= 24'h7f007f;
		12'd1995: rd_data_1 <= 24'h7f007f;
		12'd1996: rd_data_1 <= 24'h7f007f;
		12'd1997: rd_data_1 <= 24'h7f007f;
		12'd1998: rd_data_1 <= 24'h7f007f;
		12'd1999: rd_data_1 <= 24'h7f007f;
		12'd2000: rd_data_1 <= 24'h810180;
		12'd2001: rd_data_1 <= 24'h810180;
		12'd2002: rd_data_1 <= 24'h810180;
		12'd2003: rd_data_1 <= 24'h810180;
		12'd2004: rd_data_1 <= 24'h810180;
		12'd2005: rd_data_1 <= 24'h810180;
		12'd2006: rd_data_1 <= 24'h810180;
		12'd2007: rd_data_1 <= 24'h810180;
		12'd2008: rd_data_1 <= 24'h810180;
		12'd2009: rd_data_1 <= 24'h810180;
		12'd2010: rd_data_1 <= 24'h810180;
		12'd2011: rd_data_1 <= 24'h810180;
		12'd2012: rd_data_1 <= 24'h810180;
		12'd2013: rd_data_1 <= 24'h810180;
		12'd2014: rd_data_1 <= 24'h810180;
		12'd2015: rd_data_1 <= 24'h810180;
		12'd2016: rd_data_1 <= 24'h810180;
		12'd2017: rd_data_1 <= 24'h810180;
		12'd2018: rd_data_1 <= 24'h810180;
		12'd2019: rd_data_1 <= 24'h810180;
		12'd2020: rd_data_1 <= 24'h810180;
		12'd2021: rd_data_1 <= 24'h810180;
		12'd2022: rd_data_1 <= 24'h810180;
		12'd2023: rd_data_1 <= 24'h810180;
		12'd2024: rd_data_1 <= 24'h810180;
		12'd2025: rd_data_1 <= 24'h810180;
		12'd2026: rd_data_1 <= 24'h810180;
		12'd2027: rd_data_1 <= 24'h810180;
		12'd2028: rd_data_1 <= 24'h810180;
		12'd2029: rd_data_1 <= 24'h810180;
		12'd2030: rd_data_1 <= 24'h810180;
		12'd2031: rd_data_1 <= 24'h810180;
		12'd2032: rd_data_1 <= 24'h810180;
		12'd2033: rd_data_1 <= 24'h7f007f;
		12'd2034: rd_data_1 <= 24'h7f007f;
		12'd2035: rd_data_1 <= 24'h7f007f;
		12'd2036: rd_data_1 <= 24'h7f007f;
		12'd2037: rd_data_1 <= 24'h7f007f;
		12'd2038: rd_data_1 <= 24'h7f007f;
		12'd2039: rd_data_1 <= 24'h7f007f;
		12'd2040: rd_data_1 <= 24'h7f007f;
		12'd2041: rd_data_1 <= 24'h7f007f;
		12'd2042: rd_data_1 <= 24'h7f007f;
		12'd2043: rd_data_1 <= 24'h7f007f;
		12'd2044: rd_data_1 <= 24'h7f007f;
		12'd2045: rd_data_1 <= 24'h7f007f;
		12'd2046: rd_data_1 <= 24'h7f007f;
		12'd2047: rd_data_1 <= 24'h7f007f;

        endcase
    end    
        assign o_rd_data[0][2] = rd_data_0[3*bpp_p-1-:8];
        assign o_rd_data[0][1] = rd_data_0[2*bpp_p-1-:8];
        assign o_rd_data[0][0] = rd_data_0[bpp_p-1-:8];

        assign o_rd_data[1][2] = rd_data_1[3*bpp_p-1-:8];
        assign o_rd_data[1][1] = rd_data_1[2*bpp_p-1-:8];
        assign o_rd_data[1][0] = rd_data_1[bpp_p-1-:8];
endmodule