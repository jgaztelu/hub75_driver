module test_bars #(
	parameter hpixel_p = 65,
    parameter vpixel_p = 65,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

// Clock and reset
        input logic clk,
        input logic rst_n,

        /* Pixel read interface */
        input logic [addr_width_p-1:0] i_rd_addr,
        output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
        );

localparam [frame_size_p-1:0][3*bpp_p-1:0] test_bars_buf = {
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'h0000ff,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff0000,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'hff00ff,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ff00,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'h00ffff,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffff00,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff
};

    always_ff @(posedge clk) begin
        o_rd_data[0][2] <= test_bars_buf[i_rd_addr][3*bpp_p-1-:8];
        o_rd_data[0][1] <= test_bars_buf[i_rd_addr][2*bpp_p-1-:8];
        o_rd_data[0][0] <= test_bars_buf[i_rd_addr][1*bpp_p-1-:8];

        o_rd_data[1][2] <= test_bars_buf[i_rd_addr+frame_size_p/2][3*bpp_p-1-:8];
        o_rd_data[1][1] <= test_bars_buf[i_rd_addr+frame_size_p/2][2*bpp_p-1-:8];
        o_rd_data[1][0] <= test_bars_buf[i_rd_addr+frame_size_p/2][1*bpp_p-1-:8];
    end
endmodule