module shroom_rom #(
	parameter hpixel_p = 65,
    parameter vpixel_p = 65,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

// Clock and reset
        input logic clk,
        input logic rst_n,

        /* Pixel read interface */
        input logic [addr_width_p-1:0] i_rd_addr,
        output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
        );

localparam [frame_size_p-1:0][3*bpp_p-1:0] shroom_rom_buf = {
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h2ccdf1,
24'h2ccdf1,
24'h20bde9,
24'h055cae,
24'h055cae,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0668b9,
24'h0668b9,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h20bde9,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h2ccdf1,
24'h2ccdf1,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h20bde9,
24'h054fa3,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h2ccdf1,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h20bde9,
24'h054fa3,
24'h054fa3,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0668b9,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h37dbf8,
24'h2ccdf1,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h20bde9,
24'h20bde9,
24'h054fa3,
24'h054fa3,
24'h054fa3,
24'h054fa3,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0668b9,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0675c4,
24'h37dbf8,
24'h37dbf8,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h054fa3,
24'h054fa3,
24'h054fa3,
24'h054fa3,
24'h15abe2,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0668b9,
24'h0675c4,
24'h0675c4,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h37dbf8,
24'h37dbf8,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h15abe2,
24'h054fa3,
24'h054fa3,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h2ccdf1,
24'h0675c4,
24'h0675c4,
24'h0675c4,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h2ccdf1,
24'h0668b9,
24'h2ccdf1,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h2ccdf1,
24'h37dbf8,
24'h0675c4,
24'h0675c4,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h0782cf,
24'h42ecff,
24'h42ecff,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h055cae,
24'h055cae,
24'h054fa3,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h054fa3,
24'h044498,
24'h044498,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0668b9,
24'h0668b9,
24'h2ccdf1,
24'h37dbf8,
24'h37dbf8,
24'h0675c4,
24'h0675c4,
24'h0782cf,
24'h42ecff,
24'h42ecff,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h2ccdf1,
24'h2ccdf1,
24'h0668b9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h054fa3,
24'h15abe2,
24'h15abe2,
24'h054fa3,
24'h054fa3,
24'h044498,
24'h044498,
24'h044498,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h0668b9,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h055cae,
24'h054fa3,
24'h15abe2,
24'h15abe2,
24'h054fa3,
24'h054fa3,
24'h054fa3,
24'h044498,
24'h044498,
24'h044498,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h37dbf8,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h054fa3,
24'h054fa3,
24'h044498,
24'h044498,
24'h044498,
24'h044498,
24'h044498,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h20bde9,
24'h20bde9,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h054fa3,
24'h054fa3,
24'h044498,
24'h044498,
24'h044498,
24'h044498,
24'h044498,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h20bde9,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h054fa3,
24'h044498,
24'h044498,
24'h044498,
24'h044498,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h0668b9,
24'h0668b9,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h044498,
24'h044498,
24'h044498,
24'h0a9cdb,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h2ccdf1,
24'h2ccdf1,
24'h2ccdf1,
24'h0668b9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h054fa3,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h054fa3,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h055cae,
24'h054fa3,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h20bde9,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h7da9ca,
24'h7da9ca,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h15abe2,
24'h15abe2,
24'h15abe2,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h0a9cdb,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h8fb5d2,
24'h8fb5d2,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h7da9ca,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h8fb5d2,
24'h8fb5d2,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h000000,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h8fb5d2,
24'h000000,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h7da9ca,
24'h7da9ca,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h8fb5d2,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h000000,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h000000,
24'ha2c2da,
24'ha2c2da,
24'h8fb5d2,
24'h8fb5d2,
24'h7da9ca,
24'h7da9ca,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'h000000,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'ha2c2da,
24'h000000,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h8fb5d2,
24'h8fb5d2,
24'h7da9ca,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'ha2c2da,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'h000000,
24'hb4cee1,
24'h000000,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h8fb5d2,
24'h8fb5d2,
24'h8fb5d2,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'h000000,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h8fb5d2,
24'h8fb5d2,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'ha2c2da,
24'h8fb5d2,
24'h8fb5d2,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'ha2c2da,
24'h8fb5d2,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hb4cee1,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'ha2c2da,
24'ha2c2da,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'ha2c2da,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hc7dbe9,
24'hc7dbe9,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hb4cee1,
24'hb4cee1,
24'hb4cee1,
24'ha2c2da,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hc7dbe9,
24'hc7dbe9,
24'hc7dbe9,
24'hb4cee1,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'hd9e8f1,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
};

    always_ff @(posedge clk) begin
        o_rd_data[0][2] <= bulbasaur_rom_buf[i_rd_addr][3*bpp_p-1-:8];
        o_rd_data[0][1] <= bulbasaur_rom_buf[i_rd_addr][2*bpp_p-1-:8];
        o_rd_data[0][0] <= bulbasaur_rom_buf[i_rd_addr][1*bpp_p-1-:8];

        o_rd_data[1][2] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][3*bpp_p-1-:8];
        o_rd_data[1][1] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][2*bpp_p-1-:8];
        o_rd_data[1][0] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][1*bpp_p-1-:8];
    end
endmodule