module bulbasaur_rom #(
	parameter hpixel_p = 64,
    parameter vpixel_p = 64,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

// Clock and reset
        input logic clk,
        input logic rst_n,

        /* Pixel read interface */
        input logic [addr_width_p-1:0] i_rd_addr,
        output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
        );

localparam [frame_size_p-1:0][3*bpp_p-1:0] bulbasaur_rom_buf = {
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8126847,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8126847,
24'd8126847,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454269,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8257665,
24'd8126847,
24'd8126847,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8454271,
24'd8585343,
24'd8454273,
24'd8454273,
24'd8454271,
24'd8323197,
24'd8257917,
24'd8192125,
24'd8585603,
24'd8585345,
24'd8323201,
24'd8257663,
24'd8257663,
24'd8257917,
24'd8257917,
24'd8257915,
24'd8257915,
24'd8127097,
24'd7931253,
24'd8062071,
24'd8323195,
24'd8454271,
24'd8323201,
24'd8257665,
24'd8126847,
24'd8126847,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8126847,
24'd7799935,
24'd7930749,
24'd8585341,
24'd8585341,
24'd8127101,
24'd8127101,
24'd8650877,
24'd8847489,
24'd8781959,
24'd8650885,
24'd8585343,
24'd8323195,
24'd8522368,
24'd7798902,
24'd9044104,
24'd9109641,
24'd8980620,
24'd8389765,
24'd8192894,
24'd8061306,
24'd7864434,
24'd7995761,
24'd8390772,
24'd7603303,
24'd7542378,
24'd7080291,
24'd8192626,
24'd8257656,
24'd8257669,
24'd8061317,
24'd8061569,
24'd8126847,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd7930751,
24'd8061567,
24'd8650879,
24'd8650879,
24'd8061567,
24'd8061567,
24'd8585343,
24'd8781955,
24'd8781959,
24'd8650887,
24'd8454273,
24'd8061051,
24'd7667828,
24'd7733365,
24'd8586115,
24'd7995517,
24'd7473530,
24'd6292074,
24'd6489449,
24'd7542389,
24'd6753123,
24'd7674477,
24'd7279973,
24'd6427990,
24'd5645644,
24'd6961250,
24'd6623838,
24'd6619233,
24'd7538042,
24'd7799935,
24'd8061821,
24'd8127101,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257665,
24'd8257665,
24'd8323201,
24'd8323201,
24'd8323201,
24'd8323201,
24'd8257665,
24'd8323201,
24'd8650883,
24'd8585347,
24'd8061315,
24'd7931012,
24'd8126597,
24'd8323205,
24'd8585349,
24'd8454277,
24'd8126599,
24'd8323719,
24'd8651910,
24'd8259198,
24'd6817133,
24'd6493549,
24'd5841513,
24'd4923741,
24'd4726870,
24'd4924245,
24'd4463944,
24'd5122126,
24'd4595780,
24'd5850966,
24'd4017977,
24'd9348237,
24'd985362,
24'd2687020,
24'd6295388,
24'd7604591,
24'd7931253,
24'd8127097,
24'd8257917,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257665,
24'd8257665,
24'd8323201,
24'd8323201,
24'd8323201,
24'd8323201,
24'd8257665,
24'd8323201,
24'd8323203,
24'd8323203,
24'd7864449,
24'd7996292,
24'd8061317,
24'd8126851,
24'd8323201,
24'd8323201,
24'd8061315,
24'd7734655,
24'd7670904,
24'd6557540,
24'd5382232,
24'd7889025,
24'd7631237,
24'd7962250,
24'd6909558,
24'd4738897,
24'd4870733,
24'd4673350,
24'd4739397,
24'd9414795,
24'd5342795,
24'd5409617,
24'd3824705,
24'd7432822,
24'd4852806,
24'd7211878,
24'd7668595,
24'd8127101,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd7733370,
24'd8391815,
24'd7274615,
24'd7996544,
24'd7864442,
24'd8389505,
24'd7471221,
24'd8324225,
24'd8783748,
24'd8915329,
24'd8456314,
24'd7080807,
24'd5710681,
24'd7825785,
24'd6912612,
24'd10865827,
24'd10801579,
24'd10407334,
24'd10210208,
24'd10407582,
24'd10934432,
24'd8829309,
24'd8171376,
24'd8698487,
24'd5146949,
24'd8303996,
24'd3825983,
24'd6975343,
24'd2949165,
24'd7411571,
24'd7405690,
24'd8652943,
24'd8323458,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd7799933,
24'd7608195,
24'd6559356,
24'd5770609,
24'd6886524,
24'd7276149,
24'd7932538,
24'd7801209,
24'd8064638,
24'd7998843,
24'd7802997,
24'd7148135,
24'd5511505,
24'd7761791,
24'd11521722,
24'd10804394,
24'd10018207,
24'd9952932,
24'd9755553,
24'd9689755,
24'd9821850,
24'd9427088,
24'd10348442,
24'd4361531,
24'd4887107,
24'd8505216,
24'd8371842,
24'd5473114,
24'd4740941,
24'd1966113,
24'd6033504,
24'd7603583,
24'd8257673,
24'd8454276,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8323197,
24'd7211641,
24'd4463210,
24'd3746156,
24'd4339062,
24'd4400749,
24'd6168434,
24'd6361963,
24'd6625134,
24'd6032998,
24'd5967972,
24'd5050711,
24'd5321567,
24'd7500165,
24'd11257794,
24'd10078901,
24'd9491379,
24'd9559221,
24'd9624242,
24'd1004843,
24'd12546,
24'd3768653,
24'd4690005,
24'd4427085,
24'd9822109,
24'd7586685,
24'd6601332,
24'd6929019,
24'd5278297,
24'd4086339,
24'd1313307,
24'd5775708,
24'd7933050,
24'd9045384,
24'd8519808,
24'd8454528,
24'd8519810,
24'd8519810,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8323197,
24'd6753909,
24'd8024491,
24'd11653874,
24'd11194861,
24'd3230058,
24'd4011104,
24'd4862050,
24'd7033478,
24'd7034248,
24'd6574464,
24'd6117757,
24'd4744303,
24'd4157545,
24'd4029802,
24'd2585176,
24'd2454620,
24'd152119,
24'd875324,
24'd10019520,
24'd9293485,
24'd11526,
24'd9030812,
24'd9361310,
24'd9230744,
24'd9100952,
24'd6932866,
24'd6404984,
24'd7518591,
24'd3499069,
24'd6782324,
24'd2100009,
24'd6426976,
24'd7602288,
24'd8454526,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8323197,
24'd8454269,
24'd6557809,
24'd6977433,
24'd10610149,
24'd9232080,
24'd9955287,
24'd3765099,
24'd3630949,
24'd10605272,
24'd10672348,
24'd10279128,
24'd10017748,
24'd9890264,
24'd7590841,
24'd6934706,
24'd7066292,
24'd22589,
24'd9694416,
24'd9694666,
24'd10217415,
24'd10143924,
24'd8203,
24'd10343597,
24'd9557406,
24'd9297298,
24'd8707469,
24'd6865785,
24'd6602618,
24'd7258235,
24'd2716472,
24'd4752734,
24'd6323573,
24'd2229033,
24'd6953834,
24'd8061819,
24'd8716422,
24'd8650884,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8454269,
24'd6361711,
24'd6849177,
24'd9167568,
24'd3776894,
24'd8119997,
24'd9234628,
24'd9628621,
24'd8708814,
24'd8643793,
24'd3577214,
24'd3709311,
24'd3316606,
24'd8581843,
24'd6150582,
24'd5886640,
24'd7724738,
24'd8512454,
24'd8710853,
24'd7654315,
24'd9422002,
24'd8205,
24'd10934199,
24'd9621918,
24'd9692054,
24'd9431187,
24'd7259000,
24'd7324542,
24'd7061622,
24'd3245376,
24'd1468465,
24'd5738609,
24'd1252130,
24'd5054034,
24'd7538805,
24'd8650884,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8257915,
24'd8323195,
24'd8323195,
24'd8323195,
24'd8127099,
24'd5969517,
24'd6391193,
24'd1997414,
24'd8579783,
24'd9171915,
24'd9235399,
24'd8840902,
24'd8383698,
24'd3449226,
24'd4431753,
24'd3970173,
24'd4365701,
24'd8580046,
24'd7599311,
24'd5691828,
24'd6937275,
24'd6738354,
24'd7134649,
24'd6672301,
24'd7194028,
24'd5018234,
24'd9481,
24'd10014625,
24'd9757338,
24'd9298834,
24'd7783035,
24'd8111232,
24'd7060341,
24'd4165967,
24'd1600819,
24'd5083498,
24'd5666409,
24'd1771814,
24'd6754409,
24'd8192892,
24'd8454528,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8519810,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8127099,
24'd8257915,
24'd8454267,
24'd8257915,
24'd7800187,
24'd5511533,
24'd4747395,
24'd8512205,
24'd8251332,
24'd7856055,
24'd9366215,
24'd9235147,
24'd3711882,
24'd2725246,
24'd3971715,
24'd3378806,
24'd8642246,
24'd9040084,
24'd7927763,
24'd6480317,
24'd6014633,
24'd7131317,
24'd6805686,
24'd6477237,
24'd6739128,
24'd3641206,
24'd7942,
24'd10737069,
24'd9362328,
24'd7981952,
24'd8044665,
24'd8438911,
24'd7520378,
24'd4100173,
24'd3968596,
24'd1729588,
24'd5080162,
24'd659990,
24'd6035549,
24'd7800948,
24'd8127099,
24'd8454528,
24'd8585347,
24'd8585347,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8127101,
24'd8061819,
24'd8127099,
24'd8323193,
24'd8192122,
24'd7473532,
24'd4856169,
24'd4024441,
24'd8380618,
24'd8384200,
24'd9041099,
24'd9826252,
24'd8837822,
24'd4102020,
24'd3774341,
24'd3842183,
24'd8711633,
24'd8580046,
24'd8843988,
24'd8647636,
24'd7264187,
24'd4824455,
24'd4034169,
24'd6998963,
24'd6278323,
24'd6740673,
24'd3841413,
24'd8460,
24'd10933428,
24'd7519104,
24'd7455096,
24'd8175994,
24'd8241787,
24'd5152089,
24'd4232275,
24'd4033874,
24'd2125366,
24'd4493142,
24'd6588015,
24'd3080239,
24'd7212393,
24'd7800437,
24'd8126588,
24'd8585347,
24'd8585347,
24'd8323199,
24'd8257917,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8127101,
24'd8061819,
24'd8127099,
24'd8061045,
24'd8324221,
24'd6818169,
24'd7356817,
24'd3163483,
24'd10018768,
24'd6933418,
24'd8316606,
24'd8905664,
24'd9233352,
24'd9429713,
24'd9496279,
24'd7987142,
24'd8712659,
24'd8120779,
24'd7262390,
24'd10151122,
24'd4289898,
24'd12047826,
24'd11786453,
24'd1070668,
24'd7458751,
24'd3383181,
24'd3906697,
24'd5343354,
24'd9739,
24'd7452546,
24'd7389049,
24'd7585138,
24'd4230978,
24'd4365140,
24'd3443532,
24'd4362324,
24'd2059053,
24'd4627283,
24'd5078356,
24'd2557219,
24'd6754913,
24'd7669362,
24'd7995516,
24'd8585348,
24'd8585348,
24'd8192124,
24'd8061306,
24'd8257917,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8127101,
24'd7930749,
24'd8061821,
24'd8650876,
24'd8127612,
24'd6556537,
24'd5841009,
24'd6902132,
24'd7373443,
24'd9689537,
24'd7722672,
24'd9368013,
24'd8840906,
24'd9299156,
24'd4430220,
24'd3577984,
24'd8316105,
24'd6671536,
24'd10281938,
24'd5331295,
24'd7557734,
24'd6105409,
24'd16773119,
24'd12310495,
24'd1070418,
24'd4101005,
24'd3310458,
24'd5409408,
24'd7174,
24'd1727789,
24'd5020249,
24'd4035139,
24'd4497743,
24'd3512398,
24'd3050313,
24'd4887898,
24'd2321194,
24'd4034878,
24'd5539922,
24'd2165273,
24'd6493531,
24'd7407728,
24'd7995516,
24'd8585350,
24'd8585348,
24'd8192124,
24'd8061306,
24'd8257917,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8257917,
24'd8127101,
24'd8061821,
24'd8127101,
24'd8126582,
24'd7538294,
24'd5838960,
24'd5646696,
24'd8079211,
24'd9205889,
24'd11132618,
24'd7590319,
24'd8580296,
24'd8776655,
24'd3904646,
24'd3509118,
24'd3314040,
24'd8841419,
24'd7064497,
24'd11263189,
24'd7951979,
24'd9911650,
24'd8655932,
24'd16769791,
24'd16645631,
24'd1461331,
24'd4822677,
24'd3968906,
24'd4490623,
24'd11035,
24'd1004082,
24'd4362589,
24'd3838539,
24'd3576905,
24'd3182411,
24'd4167511,
24'd2584884,
24'd4361031,
24'd4560452,
24'd5407055,
24'd2492191,
24'd6689633,
24'd7538546,
24'd7995516,
24'd8585348,
24'd8585348,
24'd8192124,
24'd8061306,
24'd8257917,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8126847,
24'd8061567,
24'd8126847,
24'd8257917,
24'd8061049,
24'd6753389,
24'd7033984,
24'd13878235,
24'd9194857,
24'd16772604,
24'd6195578,
24'd8774596,
24'd8843986,
24'd8777943,
24'd4364429,
24'd4363914,
24'd8381636,
24'd9171150,
24'd9233102,
24'd6916235,
24'd8734567,
24'd16766207,
24'd9766450,
24'd8591161,
24'd16775167,
24'd11262691,
24'd3641742,
24'd4170394,
24'd4231562,
24'd807241,
24'd4294525,
24'd743486,
24'd3641180,
24'd3904087,
24'd3967570,
24'd5347938,
24'd1795883,
24'd4229706,
24'd5084752,
24'd6060124,
24'd3604533,
24'd7406703,
24'd8523138,
24'd7929976,
24'd8323201,
24'd8323201,
24'd8257917,
24'd8127101,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8061567,
24'd8061567,
24'd8126847,
24'd8257663,
24'd8061308,
24'd6097510,
24'd5921397,
24'd16121599,
24'd5973049,
24'd16772604,
24'd5868410,
24'd7461048,
24'd8187598,
24'd8515800,
24'd8708564,
24'd8906197,
24'd9107156,
24'd8382663,
24'd7851708,
24'd6390661,
24'd6105411,
24'd16769279,
24'd15890839,
24'd13596045,
24'd16774399,
24'd11591400,
24'd4167316,
24'd2986889,
24'd4233874,
24'd2783862,
24'd4952980,
24'd4492935,
24'd21305,
24'd4363632,
24'd4360804,
24'd2189372,
24'd3901773,
24'd4821330,
24'd5079119,
24'd1052688,
24'd6360929,
24'd8324223,
24'd8456064,
24'd8192894,
24'd8257663,
24'd8257663,
24'd8127101,
24'd8127101,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8126849,
24'd8061569,
24'd8061567,
24'd8061567,
24'd8061048,
24'd7018614,
24'd5922433,
24'd10664128,
24'd5057852,
24'd4009523,
24'd4427640,
24'd6215860,
24'd6084535,
24'd5952183,
24'd6805697,
24'd6542526,
24'd5755059,
24'd6214326,
24'd6868408,
24'd5410440,
24'd3617852,
24'd5911099,
24'd11962760,
24'd10980490,
24'd12570840,
24'd5670799,
24'd5216409,
24'd4298900,
24'd3906195,
24'd3904655,
24'd4492429,
24'd4820880,
24'd4493968,
24'd284496,
24'd350025,
24'd3968878,
24'd4956514,
24'd5214291,
24'd6254685,
24'd2754341,
24'd7608180,
24'd8390017,
24'd8324223,
24'd8455810,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323201,
24'd8257667,
24'd8126851,
24'd7930751,
24'd8061567,
24'd8520321,
24'd7082872,
24'd3748707,
24'd5672,
24'd11577782,
24'd10857646,
24'd9094584,
24'd7458999,
24'd6607799,
24'd6412475,
24'd6148535,
24'd6410938,
24'd6280122,
24'd6870975,
24'd7328444,
24'd8505529,
24'd10138797,
24'd11515823,
24'd10332567,
24'd10006432,
24'd6062723,
24'd5934998,
24'd938580,
24'd4033931,
24'd3642253,
24'd3904655,
24'd5085335,
24'd5084055,
24'd4689814,
24'd4953500,
24'd4757654,
24'd612677,
24'd4296794,
24'd5867358,
24'd1640473,
24'd6693476,
24'd7210092,
24'd8192894,
24'd8455810,
24'd8192894,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323201,
24'd8323205,
24'd8257669,
24'd7930751,
24'd8061821,
24'd8126588,
24'd7015030,
24'd4794219,
24'd7436187,
24'd4896,
24'd2767681,
24'd11645372,
24'd11321538,
24'd4757123,
24'd6869942,
24'd7789762,
24'd1802086,
24'd6473389,
24'd7787451,
24'd7652269,
24'd8569003,
24'd9156004,
24'd10536885,
24'd3763289,
24'd1001530,
24'd8480,
24'd7457,
24'd4558478,
24'd3902345,
24'd2389106,
24'd4494482,
24'd4231310,
24'd4229511,
24'd1134415,
24'd1396817,
24'd5214610,
24'd4754563,
24'd1396787,
24'd531223,
24'd5710433,
24'd6948719,
24'd7931001,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8585351,
24'd8454279,
24'd8126847,
24'd8061821,
24'd8323712,
24'd7735934,
24'd5180003,
24'd4598373,
24'd7306132,
24'd15728639,
24'd3680572,
24'd3617600,
24'd9419956,
24'd9225654,
24'd10009524,
24'd10664887,
24'd10138797,
24'd5729637,
24'd3819326,
24'd1056274,
24'd136969,
24'd6926,
24'd13762559,
24'd2650218,
24'd5279374,
24'd5344142,
24'd5083539,
24'd4690064,
24'd743767,
24'd4033931,
24'd4692372,
24'd4690830,
24'd1726034,
24'd1593934,
24'd1266514,
24'd5477520,
24'd5211513,
24'd3095882,
24'd5906795,
24'd6619502,
24'd7931003,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454275,
24'd8650889,
24'd8650887,
24'd8454271,
24'd8257915,
24'd7733372,
24'd8325509,
24'd7932538,
24'd6558313,
24'd4861018,
24'd7961746,
24'd7176332,
24'd5268584,
24'd3159610,
24'd4532278,
24'd7347772,
24'd9117506,
24'd7934253,
24'd8329520,
24'd8133163,
24'd7217451,
24'd5451059,
24'd3619907,
24'd3960697,
24'd4295059,
24'd4688529,
24'd5477016,
24'd5869207,
24'd936783,
24'd4100494,
24'd4102289,
24'd4034953,
24'd5414807,
24'd4755591,
24'd1070670,
24'd545356,
24'd4492168,
24'd5214092,
24'd6324366,
24'd5059172,
24'd6165863,
24'd7538805,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8650887,
24'd8650885,
24'd8585341,
24'd8323197,
24'd7471225,
24'd7864444,
24'd8650876,
24'd7799663,
24'd6955628,
24'd2360630,
24'd856883,
24'd7306898,
24'd7762305,
24'd7753312,
24'd7082547,
24'd11681635,
24'd14970770,
24'd14971533,
24'd14249345,
24'd13137794,
24'd8542816,
24'd7698560,
24'd5538961,
24'd4491929,
24'd5544356,
24'd8747,
24'd10548,
24'd4819086,
24'd3706761,
24'd4168849,
24'd4034181,
24'd4427910,
24'd2717806,
24'd4494216,
24'd4625034,
24'd4690316,
24'd5018516,
24'd5538961,
24'd3422296,
24'd4528470,
24'd7211891,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454273,
24'd8454273,
24'd8454269,
24'd8323197,
24'd8061056,
24'd8192128,
24'd8454270,
24'd8388730,
24'd8063352,
24'd6688366,
24'd5249644,
24'd1114167,
24'd3100,
24'd7046790,
24'd7240828,
24'd7895421,
24'd8417920,
24'd8614268,
24'd9075836,
24'd8881276,
24'd7570293,
24'd6720126,
24'd10024,
24'd9516,
24'd9009,
24'd4885142,
24'd4164754,
24'd3246214,
24'd2062192,
24'd3574659,
24'd4427140,
24'd611401,
24'd4167302,
24'd4101255,
24'd4558474,
24'd806992,
24'd4360331,
24'd4949137,
24'd6586521,
24'd1836862,
24'd6753907,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323199,
24'd8192126,
24'd8192128,
24'd8454270,
24'd8585342,
24'd7995507,
24'd8127614,
24'd6490230,
24'd5450870,
24'd6390420,
24'd10781,
24'd12317,
24'd7953,
24'd8738,
24'd9766,
24'd7958,
24'd8205,
24'd9485,
24'd7948,
24'd4754565,
24'd4886674,
24'd4426386,
24'd4165013,
24'd3510161,
24'd3445392,
24'd21582,
24'd4296072,
24'd5148298,
24'd12072,
24'd3576197,
24'd4233872,
24'd1136727,
24'd1397847,
24'd1003862,
24'd4488584,
24'd6458012,
24'd1511232,
24'd6688627,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8192126,
24'd8192126,
24'd8454270,
24'd8585342,
24'd8650878,
24'd7602293,
24'd7539838,
24'd9199275,
24'd9354442,
24'd6603440,
24'd7064758,
24'd4167302,
24'd938317,
24'd5409928,
24'd5608325,
24'd5083775,
24'd4758406,
24'd3640445,
24'd4887439,
24'd20044,
24'd7066574,
24'd6475466,
24'd3643798,
24'd3772558,
24'd4296333,
24'd1135443,
24'd5658,
24'd4949641,
24'd4168597,
24'd2919046,
24'd1004375,
24'd1067088,
24'd1199186,
24'd5473934,
24'd6062475,
24'd655658,
24'd6688625,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8192126,
24'd8192126,
24'd8454270,
24'd8454270,
24'd9046406,
24'd7929976,
24'd7997309,
24'd5512300,
24'd4222334,
24'd3446405,
24'd6737592,
24'd6932918,
24'd3967620,
24'd872270,
24'd12069,
24'd4686971,
24'd5081225,
24'd4556168,
24'd413004,
24'd4364177,
24'd3382931,
24'd6278595,
24'd7328460,
24'd3706765,
24'd4492429,
24'd1659223,
24'd6953,
24'd6130067,
24'd4627353,
24'd3971734,
24'd1071965,
24'd542285,
24'd1463127,
24'd5802386,
24'd6322567,
24'd2231609,
24'd6884975,
24'd8257917,
24'd8257917,
24'd8257917,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8454271,
24'd8585343,
24'd8519806,
24'd8257660,
24'd8324221,
24'd6035308,
24'd4614012,
24'd3642244,
24'd6473651,
24'd6999484,
24'd4231821,
24'd5083024,
24'd6460048,
24'd268580,
24'd1642038,
24'd855348,
24'd1463125,
24'd4365199,
24'd3640708,
24'd3773323,
24'd7393991,
24'd4300183,
24'd3702402,
24'd1656658,
24'd267563,
24'd6782866,
24'd4622988,
24'd4102291,
24'd4101007,
24'd613209,
24'd4756373,
24'd5342096,
24'd987951,
24'd4330575,
24'd7211889,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8454271,
24'd8585343,
24'd8650878,
24'd8519806,
24'd8454780,
24'd6558572,
24'd6977683,
24'd8833988,
24'd7391159,
24'd7590337,
24'd8049614,
24'd4426125,
24'd6390409,
24'd1445161,
24'd5380700,
24'd4662368,
24'd5737876,
24'd7260856,
24'd4362630,
24'd4231560,
24'd6670780,
24'd3640969,
24'd5736340,
24'd3425375,
24'd3221836,
24'd789543,
24'd3630183,
24'd5149321,
24'd2846827,
24'd4951437,
24'd3172980,
24'd6783132,
24'd2360632,
24'd5901916,
24'd7735157,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8454271,
24'd8585343,
24'd8716414,
24'd8650878,
24'd8454780,
24'd6885740,
24'd4140371,
24'd4877168,
24'd9226947,
24'd4495500,
24'd7130311,
24'd4690326,
24'd6518147,
24'd1900582,
24'd6100072,
24'd4988519,
24'd4947590,
24'd7524796,
24'd7324851,
24'd7852223,
24'd6408376,
24'd4756112,
24'd987438,
24'd5056342,
24'd5318235,
24'd4598864,
24'd12175300,
24'd2245171,
24'd12441300,
24'd2899017,
24'd12962282,
24'd4663905,
24'd6097760,
24'd7537258,
24'd8127097,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8454271,
24'd8585343,
24'd8716418,
24'd8716416,
24'd8454780,
24'd7277936,
24'd5646687,
24'd16709887,
24'd2835021,
24'd14942207,
24'd1265496,
24'd5931668,
24'd1837616,
24'd5511514,
24'd6886774,
24'd5052779,
24'd2575197,
24'd8177339,
24'd5148548,
24'd8832443,
24'd5149582,
24'd6588054,
24'd2228271,
24'd6362717,
24'd6164318,
24'd5509716,
24'd2294560,
24'd1771032,
24'd2295589,
24'd2424879,
24'd3080254,
24'd6100072,
24'd7932018,
24'd8782714,
24'd8454267,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8454271,
24'd8585345,
24'd8716424,
24'd8650888,
24'd8323712,
24'd7473782,
24'd6164833,
24'd3145782,
24'd1638434,
24'd2165036,
24'd1376806,
24'd2622775,
24'd6231912,
24'd6950772,
24'd6556791,
24'd6038392,
24'd16120575,
24'd2244682,
24'd15990783,
24'd3226437,
24'd16118783,
24'd2295607,
24'd6100322,
24'd7211630,
24'd7734390,
24'd7734390,
24'd7146348,
24'd6950248,
24'd7015532,
24'd7146096,
24'd7211380,
24'd7538294,
24'd8061306,
24'd8388732,
24'd8323197,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8454271,
24'd8585345,
24'd8716424,
24'd8650888,
24'd8323712,
24'd7800696,
24'd7343727,
24'd6623074,
24'd6164568,
24'd6231126,
24'd6361431,
24'd6687584,
24'd7867002,
24'd7603585,
24'd7080321,
24'd6099318,
24'd2687044,
24'd2032949,
24'd2097195,
24'd2949168,
24'd3539001,
24'd6362213,
24'd7146350,
24'd7865208,
24'd8388736,
24'd8585346,
24'd8388736,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8454271,
24'd8454271,
24'd8650880,
24'd8650880,
24'd8454780,
24'd8193144,
24'd7603055,
24'd7801200,
24'd7736942,
24'd7670382,
24'd8325496,
24'd8521857,
24'd8061058,
24'd8127112,
24'd7405698,
24'd7604100,
24'd7277436,
24'd7475579,
24'd7277686,
24'd7276919,
24'd7341429,
24'd7669112,
24'd7865210,
24'd8061308,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257660,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8454269,
24'd8650876,
24'd8520060,
24'd8520060,
24'd8454778,
24'd8718207,
24'd8258167,
24'd8061045,
24'd8323449,
24'd8126584,
24'd8716421,
24'd7995519,
24'd8389001,
24'd7995524,
24'd8323206,
24'd8061054,
24'd8061054,
24'd8192129,
24'd8783498,
24'd8061052,
24'd8389251,
24'd8192126,
24'd8192126,
24'd8192126,
24'd8192124,
24'd8257660,
24'd8257660,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8257662,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8454269,
24'd8520060,
24'd8520060,
24'd8520060,
24'd8650878,
24'd8650878,
24'd8716416,
24'd8716416,
24'd8650880,
24'd8257665,
24'd8126849,
24'd8323199,
24'd8519806,
24'd8388732,
24'd8388734,
24'd8257664,
24'd8192126,
24'd8127097,
24'd8127351,
24'd8127097,
24'd8258169,
24'd8257915,
24'd8257917,
24'd8257663,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323197,
24'd8323197,
24'd8519808,
24'd8519808,
24'd8519808,
24'd8650880,
24'd8650882,
24'd8716418,
24'd8716418,
24'd8519810,
24'd8061569,
24'd8061567,
24'd8257917,
24'd8454269,
24'd8388732,
24'd8257660,
24'd8061054,
24'd8061308,
24'd8258167,
24'd8323701,
24'd8323701,
24'd8323447,
24'd8323195,
24'd8257917,
24'd8257917,
24'd8257663,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454271,
24'd8454273,
24'd8519814,
24'd8519816,
24'd8519814,
24'd8454276,
24'd8323458,
24'd8323458,
24'd8192640,
24'd8192640,
24'd8127101,
24'd8257917,
24'd8257665,
24'd8257667,
24'd8061058,
24'd7930240,
24'd7734140,
24'd7930490,
24'd8650873,
24'd8978553,
24'd8847481,
24'd8650875,
24'd8454267,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454271,
24'd8454273,
24'd8519814,
24'd8519816,
24'd8454278,
24'd8323460,
24'd8192642,
24'd8127360,
24'd8127360,
24'd8127614,
24'd8257917,
24'd8323197,
24'd8257665,
24'd8257667,
24'd8061058,
24'd7864704,
24'd7734140,
24'd8061308,
24'd8781949,
24'd8978557,
24'd8847485,
24'd8781949,
24'd8585341,
24'd8323197,
24'd8257917,
24'd8257917,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454274,
24'd8454274,
24'd8454274,
24'd8454274,
24'd8323712,
24'd8323712,
24'd8323712,
24'd8323712,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454274,
24'd8257665,
24'd8257663,
24'd8126847,
24'd8257663,
24'd8454271,
24'd8585343,
24'd8585343,
24'd8454271,
24'd8454271,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8454528,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199,
24'd8323199};

    always_ff @(posedge clk) begin
        o_rd_data[0][2] <= bulbasaur_rom_buf[i_rd_addr][23:16];
        o_rd_data[0][1] <= bulbasaur_rom_buf[i_rd_addr][15:8];
        o_rd_data[0][0] <= bulbasaur_rom_buf[i_rd_addr][7:0];

        o_rd_data[1][2] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][23:16];
        o_rd_data[1][1] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][15:8];
        o_rd_data[1][0] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][7:0];
    end
endmodule