module bulbasaur_rom #(
    parameter hpixel_p = 64,
    parameter vpixel_p = 64,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

    // Clock and reset
    input logic clk,
    input logic rst_n,

    /* Pixel read interface */
    input logic [addr_width_p-1:0] i_rd_addr,
    output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
    );

	localparam [frame_size_p-1:0][3*bpp_p-1:0] bulbasaur_rom_buf = {
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h80007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h80007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h80007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h80007f,
		24'h81007f,
		24'h82007f,
		24'h83007f,
		24'h82007f,
		24'h7f007f,
		24'h7d017f,
		24'h7d017f,
		24'h7e0080,
		24'h7f0082,
		24'h810081,
		24'h810180,
		24'h810180,
		24'h800180,
		24'h7f0280,
		24'h7f0280,
		24'h7f0280,
		24'h800181,
		24'h810082,
		24'h810082,
		24'h810082,
		24'h810081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e017e,
		24'h7e017d,
		24'h7e007d,
		24'h81007d,
		24'h85007d,
		24'h87007d,
		24'h88007d,
		24'h88007d,
		24'h81007c,
		24'h78027c,
		24'h76027e,
		24'h790081,
		24'h7d0083,
		24'h7e0082,
		24'h7e007f,
		24'h7f007d,
		24'h7d027d,
		24'h7c047f,
		24'h7c0380,
		24'h7c0381,
		24'h7e0283,
		24'h800185,
		24'h810087,
		24'h820088,
		24'h820085,
		24'h810080,
		24'h81007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e017e,
		24'h7e017d,
		24'h7e007d,
		24'h80007c,
		24'h83007b,
		24'h86007a,
		24'h89007a,
		24'h880079,
		24'h7e0179,
		24'h77037b,
		24'h77027e,
		24'h7a0081,
		24'h7c0083,
		24'h7e0082,
		24'h7e007f,
		24'h7d017d,
		24'h7c027e,
		24'h7d0280,
		24'h7d0281,
		24'h7e0182,
		24'h800182,
		24'h810085,
		24'h820087,
		24'h820088,
		24'h820085,
		24'h810080,
		24'h81007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e017e,
		24'h7e017d,
		24'h7f007c,
		24'h7f0079,
		24'h800276,
		24'h800275,
		24'h800276,
		24'h7c027a,
		24'h7a007d,
		24'h7b007d,
		24'h7e007c,
		24'h80007d,
		24'h80007d,
		24'h7d017e,
		24'h7a0280,
		24'h7d0182,
		24'h830082,
		24'h840082,
		24'h840082,
		24'h840081,
		24'h830081,
		24'h820081,
		24'h820081,
		24'h810080,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e017e,
		24'h7e017c,
		24'h7e0279,
		24'h7d0278,
		24'h7c0377,
		24'h7c0377,
		24'h7c017c,
		24'h7d007f,
		24'h7f007f,
		24'h80007c,
		24'h81007c,
		24'h81007d,
		24'h7e0080,
		24'h7b0181,
		24'h800082,
		24'h850081,
		24'h860081,
		24'h850080,
		24'h84007e,
		24'h83007d,
		24'h82017c,
		24'h82017c,
		24'h82017c,
		24'h81007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007d,
		24'h7e007c,
		24'h7d007c,
		24'h7d007d,
		24'h7d007e,
		24'h7d007e,
		24'h7f0181,
		24'h7e017e,
		24'h810483,
		24'h820385,
		24'h7c007f,
		24'h7c007d,
		24'h7e0082,
		24'h7e0084,
		24'h7e0086,
		24'h7e0184,
		24'h7e0081,
		24'h810081,
		24'h7e0079,
		24'h7f007a,
		24'h7d0077,
		24'h81037b,
		24'h85057f,
		24'h81017a,
		24'h82017c,
		24'h83017c,
		24'h84007c,
		24'h80007d,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007c,
		24'h7e007d,
		24'h7e007d,
		24'h7e007e,
		24'h7c007d,
		24'h7a017c,
		24'h78037b,
		24'h76047a,
		24'h76077d,
		24'h770a7d,
		24'h780e7e,
		24'h770e7f,
		24'h760883,
		24'h740284,
		24'h770086,
		24'h7c0186,
		24'h7f0283,
		24'h840781,
		24'h7d0776,
		24'h780a70,
		24'h790b71,
		24'h780672,
		24'h780373,
		24'h80047a,
		24'h82017c,
		24'h84007f,
		24'h83007f,
		24'h81007f,
		24'h81007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007e,
		24'h7e007e,
		24'h7f007e,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h800080,
		24'h820082,
		24'h820081,
		24'h7d007d,
		24'h740574,
		24'h6e1170,
		24'h49004c,
		24'h330036,
		24'h2a0030,
		24'h240033,
		24'h27003e,
		24'h41005b,
		24'h6a0d80,
		24'h710583,
		24'h790581,
		24'h760875,
		24'h6d0d64,
		24'h69125e,
		24'h66135d,
		24'h681062,
		24'h6e0e6a,
		24'h740a72,
		24'h7a057b,
		24'h810182,
		24'h850088,
		24'h850086,
		24'h830080,
		24'h81007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007c,
		24'h7d007c,
		24'h780379,
		24'h75077a,
		24'h750978,
		24'h740975,
		24'h730b72,
		24'h740a73,
		24'h790479,
		24'h7b027b,
		24'h750575,
		24'h6c116e,
		24'h34003f,
		24'h9980a2,
		24'h797283,
		24'h878691,
		24'h75818d,
		24'h76818e,
		24'had8ebe,
		24'h570a71,
		24'h6a0979,
		24'h6f1177,
		24'h520d59,
		24'h26002f,
		24'h1f0027,
		24'h1f0025,
		24'h240029,
		24'h3c0040,
		24'h6b106d,
		24'h77077b,
		24'h810183,
		24'h85008a,
		24'h850087,
		24'h830080,
		24'h81007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h80007b,
		24'h86027c,
		24'h800577,
		24'h6b1070,
		24'h3c0048,
		24'h31003a,
		24'h29002b,
		24'h280225,
		24'h24001f,
		24'h490647,
		24'h620c63,
		24'h691165,
		24'h410343,
		24'h423d60,
		24'h68939b,
		24'h76ada7,
		24'h74a9a0,
		24'h6faea4,
		24'h5e9494,
		24'h4e4473,
		24'h5b1273,
		24'h681671,
		24'h410c4a,
		24'h352e52,
		24'h315569,
		24'h51737e,
		24'h94a1ab,
		24'h565a69,
		24'hc6abc6,
		24'h55115b,
		24'h760875,
		24'h83017f,
		24'h850083,
		24'h850083,
		24'h83007f,
		24'h81007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7e017b,
		24'h7b0072,
		24'h6d0769,
		24'h481258,
		24'h9f8ebc,
		24'h44455e,
		24'h879198,
		24'h40534b,
		24'h77837d,
		24'h6d5873,
		24'h4e1e55,
		24'h59235c,
		24'h230631,
		24'h305463,
		24'h56afa6,
		24'h70cdbd,
		24'h74c7b6,
		24'h71cbb7,
		24'h5ba89f,
		24'h40416c,
		24'h59146c,
		24'h48084e,
		24'h362544,
		24'h527683,
		24'h50a2a5,
		24'h5db5ae,
		24'h6fb1a9,
		24'h7ba6a5,
		24'h606978,
		24'h481a54,
		24'h730b73,
		24'h83007e,
		24'h84007e,
		24'h85007f,
		24'h83007f,
		24'h81007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h80007e,
		24'h7b0479,
		24'h680a66,
		24'h380142,
		24'h55537c,
		24'h5a8194,
		24'h4b8086,
		24'h4d8885,
		24'h478479,
		24'h578681,
		24'h283042,
		24'h2a193f,
		24'h3c3459,
		24'h445a71,
		24'h3d7f83,
		24'h52b5a9,
		24'h59b6aa,
		24'h4a998e,
		24'h62bbaa,
		24'h6ab9b0,
		24'h51597c,
		24'h541963,
		24'h390b42,
		24'h34384c,
		24'h59898f,
		24'h58aaab,
		24'h78d6cd,
		24'h6ac4b4,
		24'h7cc8bc,
		24'h729fa5,
		24'h604b7b,
		24'h6d086e,
		24'h83007e,
		24'h83007e,
		24'h84007e,
		24'h83007f,
		24'h81007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h80007e,
		24'h760776,
		24'h55135c,
		24'h13022a,
		24'h46677c,
		24'h4c8f95,
		24'h217170,
		24'h2e807c,
		24'h419891,
		24'h3f8787,
		24'h4f6f7d,
		24'h252f48,
		24'h132e41,
		24'h346c76,
		24'h3f908f,
		24'h5dbfb5,
		24'h52aea4,
		24'h33867e,
		24'h459d91,
		24'h3d8c84,
		24'h1c344d,
		24'h1d0337,
		24'h110327,
		24'h2c474e,
		24'h669d9d,
		24'h4c9696,
		24'h5ab4ab,
		24'h6ed2be,
		24'h5cbdaa,
		24'h4b9490,
		24'h53517b,
		24'h680a6e,
		24'h82017e,
		24'h80007d,
		24'h83007d,
		24'h83007f,
		24'h81007f,
		24'h7f007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7e017d,
		24'h7e017d,
		24'h7f007e,
		24'h720b75,
		24'h350a45,
		24'h424a61,
		24'h57838e,
		24'h337176,
		24'h0a4d52,
		24'h135e5f,
		24'h338e8b,
		24'h439c99,
		24'h63979f,
		24'h223d4d,
		24'h08313c,
		24'h327377,
		24'h3b8c8b,
		24'h5dbcb6,
		24'h68cfc6,
		24'h3ea69c,
		24'h3d9b92,
		24'h24716c,
		24'h164f56,
		24'h3d6775,
		24'h3c696e,
		24'h26574f,
		24'h134742,
		24'h256d6c,
		24'h52a89e,
		24'h6fd5c0,
		24'h52bba5,
		24'h2d827a,
		24'h404c71,
		24'h5f0c6c,
		24'h7e037e,
		24'h7e027c,
		24'h880684,
		24'h81007d,
		24'h80007e,
		24'h7e007e,
		24'h7d007e,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7e017d,
		24'h7e017d,
		24'h80007e,
		24'h710d77,
		24'h1a0132,
		24'h4d6676,
		24'h5f8e96,
		24'h225b61,
		24'h0d444c,
		24'h0b4b50,
		24'h247c7a,
		24'h3b9b96,
		24'h569c9f,
		24'h1a363e,
		24'h002c30,
		24'h347b7b,
		24'h419291,
		24'h3e9c98,
		24'h59c3be,
		24'h68d8d1,
		24'h32908a,
		24'h1c6664,
		24'h3d8b85,
		24'h489e90,
		24'h54a190,
		24'h4c8d7d,
		24'h427d74,
		24'h327270,
		24'h2a7a71,
		24'h60c2af,
		24'h6cd5bf,
		24'h65bcb1,
		24'h7f91b3,
		24'h7e3793,
		24'h740379,
		24'h790077,
		24'h870382,
		24'h82007e,
		24'h80007e,
		24'h7d007e,
		24'h7d007e,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7e017d,
		24'h7e017d,
		24'h80007e,
		24'h700c78,
		24'h1d053d,
		24'h4f6e83,
		24'h548893,
		24'h1a575e,
		24'h114d52,
		24'h0c4d50,
		24'h2c817c,
		24'h3d9d93,
		24'h1e5e58,
		24'h2a5856,
		24'h397976,
		24'h1c6a66,
		24'h257e7b,
		24'h359392,
		24'h3e989b,
		24'h53a9ae,
		24'h459497,
		24'h46908e,
		24'h306c5f,
		24'h093720,
		24'h0d3f28,
		24'h103c2c,
		24'h14413a,
		24'h073736,
		24'h002b24,
		24'h0f4633,
		24'h185641,
		24'h366c65,
		24'h7c8caf,
		24'h692b85,
		24'h6d0378,
		24'h7d017b,
		24'h7e0077,
		24'h83007f,
		24'h80007e,
		24'h7d007f,
		24'h7d007e,
		24'h7f007f,
		24'h7f007e,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7e017d,
		24'h7e017d,
		24'h80007e,
		24'h700c78,
		24'h210141,
		24'h576e8b,
		24'h528796,
		24'h387b82,
		24'h115356,
		24'h276c6b,
		24'h3e9087,
		24'h439d8f,
		24'h0e574b,
		24'h2e7269,
		24'h47958f,
		24'h1e746c,
		24'h1f7a75,
		24'h3a9294,
		24'h4a98a1,
		24'h2a606e,
		24'h123841,
		24'h153f41,
		24'h275148,
		24'h4b6754,
		24'h4f6251,
		24'h565e55,
		24'h535859,
		24'h4f555e,
		24'h4e585c,
		24'h495f59,
		24'h496960,
		24'h355655,
		24'h151936,
		24'h2d0550,
		24'h641478,
		24'h760977,
		24'h7e0378,
		24'h82007d,
		24'h80007f,
		24'h7d0080,
		24'h7c0080,
		24'h80007e,
		24'h80007d,
		24'h800080,
		24'h800080,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e007e,
		24'h7e017d,
		24'h7e017d,
		24'h7f007e,
		24'h730977,
		24'h3f0d51,
		24'h3d3f63,
		24'h4e798a,
		24'h4e9297,
		24'h37807d,
		24'h458f89,
		24'h4b9a8f,
		24'h36887b,
		24'h2d7c70,
		24'h39877d,
		24'h3e958b,
		24'h338e85,
		24'h408f8e,
		24'h27636b,
		24'h133842,
		24'h275762,
		24'h336c78,
		24'h2e606b,
		24'h56757a,
		24'h807d7d,
		24'h9e787a,
		24'hc7848c,
		24'hcf7b8c,
		24'hd27d96,
		24'hc3708c,
		24'h914962,
		24'h724559,
		24'h6e6370,
		24'h4f5166,
		24'h414267,
		24'h1b053a,
		24'h43054c,
		24'h781675,
		24'h7e0075,
		24'h83007e,
		24'h77007c,
		24'h75007b,
		24'h80007d,
		24'h82007e,
		24'h830084,
		24'h830085,
		24'h800080,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e017d,
		24'h7e017d,
		24'h7f017e,
		24'h750777,
		24'h5d1465,
		24'h432759,
		24'h597387,
		24'h549294,
		24'h4b938f,
		24'h28746d,
		24'h1d675e,
		24'h358076,
		24'h4e9990,
		24'h44948c,
		24'h3d968e,
		24'h429c95,
		24'h2c7374,
		24'h2b5e67,
		24'h38646c,
		24'h427f86,
		24'h4d97a2,
		24'h40828f,
		24'h45626d,
		24'h5b474f,
		24'h7f3d47,
		24'ha13b4a,
		24'ha9334a,
		24'ha72e4c,
		24'ha02348,
		24'h8b143b,
		24'h60112e,
		24'h4c3140,
		24'h4e565e,
		24'h5e757e,
		24'h4a596d,
		24'h4f3e63,
		24'h571c5e,
		24'h73096f,
		24'h81067e,
		24'h7b0481,
		24'h75007a,
		24'h80007c,
		24'h83007f,
		24'h840088,
		24'h840089,
		24'h810082,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e017d,
		24'h7e017d,
		24'h7e017d,
		24'h79057a,
		24'h68066f,
		24'h5a1d6a,
		24'h474a65,
		24'h50817d,
		24'h559791,
		24'h1b5f5c,
		24'h0b4a46,
		24'h23615b,
		24'h448b86,
		24'h499a93,
		24'h419690,
		24'h277a77,
		24'h236d6d,
		24'h46878a,
		24'h5c9b9f,
		24'h58999c,
		24'h3b8283,
		24'h71b0b4,
		24'h608182,
		24'h0b0906,
		24'h1b0e09,
		24'h361817,
		24'h523235,
		24'h71545a,
		24'h987b85,
		24'h9d838f,
		24'h828184,
		24'h708c87,
		24'h5c7373,
		24'h33323f,
		24'h6f707e,
		24'hc7d2dd,
		24'h5a4d78,
		24'h4e1361,
		24'h650770,
		24'h7d0983,
		24'h7c017f,
		24'h7c027c,
		24'h7f0080,
		24'h820088,
		24'h840087,
		24'h810081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e017d,
		24'h7e017d,
		24'h7e017d,
		24'h7c037c,
		24'h6d0073,
		24'h651c71,
		24'h1f1b30,
		24'h1d4b3a,
		24'h498a7f,
		24'h448584,
		24'h1d5858,
		24'h0a4443,
		24'h307573,
		24'h449490,
		24'h459593,
		24'h247271,
		24'h2d7c7a,
		24'h4d9b9a,
		24'h316668,
		24'h1a3d3f,
		24'h0d453e,
		24'h417e72,
		24'h719d8f,
		24'h5c7a6a,
		24'h4f7866,
		24'h548775,
		24'h609e8c,
		24'h72bca8,
		24'h68b5a2,
		24'h5daa97,
		24'h88ddc7,
		24'h73c8b1,
		24'h6d9b93,
		24'h837e8b,
		24'h817b88,
		24'h5f7478,
		24'h2b3a52,
		24'h65578b,
		24'h4e1368,
		24'h74077b,
		24'h7e017d,
		24'h7b037d,
		24'h7a0280,
		24'h7f0086,
		24'h810085,
		24'h800081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7d017d,
		24'h800480,
		24'h7e027f,
		24'h740173,
		24'h721671,
		24'h3a093d,
		24'h34453a,
		24'h2f6e43,
		24'h1d6951,
		24'h45918d,
		24'h44898e,
		24'h307379,
		24'h408588,
		24'h4a9494,
		24'h449693,
		24'h358c88,
		24'h388c88,
		24'h2b7777,
		24'h285e63,
		24'h2e5054,
		24'h436a61,
		24'h628773,
		24'h90ac9a,
		24'hb3cfc3,
		24'h98cabb,
		24'h80d2be,
		24'h72d7bf,
		24'h6ad9bf,
		24'h4fc0a6,
		24'h48b89e,
		24'h68dbbf,
		24'h5cccb0,
		24'h65bca7,
		24'h9dd3c8,
		24'h99b5b4,
		24'h6c757b,
		24'h596271,
		24'h263150,
		24'h47276a,
		24'h720a7a,
		24'h80017f,
		24'h7a027e,
		24'h79037f,
		24'h7d0184,
		24'h7e0084,
		24'h7f0081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f0481,
		24'h800581,
		24'h800481,
		24'h770d77,
		24'h4e104a,
		24'h3d313a,
		24'h538054,
		24'h51a162,
		24'h2e835d,
		24'h1e7164,
		24'h1e6e6d,
		24'h3f8c90,
		24'h4e9699,
		24'h4b9092,
		24'h409491,
		24'h399891,
		24'h3f9893,
		24'h368281,
		24'h417e83,
		24'h79a1a9,
		24'ha0adaa,
		24'hada296,
		24'h947d79,
		24'h675d5f,
		24'h618581,
		24'h68bdad,
		24'h66d4bc,
		24'h5bd1b6,
		24'h5bd2b9,
		24'h64d6bf,
		24'h5dd3b9,
		24'h5bd4b7,
		24'h60d8b8,
		24'h61ccad,
		24'h5e9283,
		24'h6c5c62,
		24'h786d7a,
		24'h4c6473,
		24'h514275,
		24'h721079,
		24'h7f007c,
		24'h7a027f,
		24'h7a037f,
		24'h7b0282,
		24'h7d0082,
		24'h7e0080,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7d017e,
		24'h7d017e,
		24'h7e007f,
		24'h7e007f,
		24'h7f0480,
		24'h80057f,
		24'h820482,
		24'h761377,
		24'h1f001d,
		24'h496248,
		24'h519055,
		24'h489858,
		24'h348254,
		24'h257053,
		24'h24745c,
		24'h1a6c5b,
		24'h3a857e,
		24'h4c9394,
		24'h3a8989,
		24'h39948d,
		24'h38988f,
		24'h3c9692,
		24'h67a7ac,
		24'hc1d9e2,
		24'hd9b7c3,
		24'hd17e8c,
		24'hce8fa2,
		24'h7b576d,
		24'h43434e,
		24'h62a89e,
		24'h70d8bf,
		24'h70e2c1,
		24'h77e5ca,
		24'h7de3d1,
		24'h78e2cf,
		24'h6ee3c7,
		24'h6be3c1,
		24'h5cc2a2,
		24'h61897d,
		24'h90707f,
		24'h674553,
		24'hcce0e5,
		24'h534871,
		24'h67086e,
		24'h7c007c,
		24'h7d017f,
		24'h7c017f,
		24'h7b0280,
		24'h7b0280,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7c027d,
		24'h7d027d,
		24'h7e0080,
		24'h7e0080,
		24'h7a017b,
		24'h820a82,
		24'h7d047c,
		24'h540653,
		24'h393539,
		24'h487f4a,
		24'h489150,
		24'h2e7a3d,
		24'h347c47,
		24'h418958,
		24'h469766,
		24'h257c50,
		24'h1b6a51,
		24'h3f8881,
		24'h2b7470,
		24'h2f807a,
		24'h3c9d93,
		24'h2d918a,
		24'h7dc1c6,
		24'hf0ffff,
		24'hd495aa,
		24'ha82744,
		24'hf19ac2,
		24'hd0a3c8,
		24'h604559,
		24'h6fa9a2,
		24'h89e8ce,
		24'h8bf4d1,
		24'h7fe1c7,
		24'h61b6ac,
		24'h6ecdbe,
		24'h88f7dc,
		24'h83f0cf,
		24'h6ec2a6,
		24'h88a29b,
		24'hf8d6eb,
		24'h89556a,
		24'hdddfeb,
		24'h59436f,
		24'h65036a,
		24'h7d007c,
		24'h7e007f,
		24'h7c017f,
		24'h7b027f,
		24'h7b027f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h800180,
		24'h800180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e017e,
		24'h7b017b,
		24'h7d007c,
		24'h810082,
		24'h820084,
		24'h7a007b,
		24'h7c097b,
		24'h720c6f,
		24'h34002f,
		24'h526750,
		24'h4f974f,
		24'h46924b,
		24'h236d2e,
		24'h408f52,
		24'h3d9254,
		24'h358f4d,
		24'h3c9655,
		24'h2b7e4d,
		24'h276f54,
		24'h0e4839,
		24'h286860,
		24'h439892,
		24'h3d9793,
		24'h468a8f,
		24'hbbd2d5,
		24'he1c2cc,
		24'h9b3657,
		24'haa3c69,
		24'hb07095,
		24'h847584,
		24'h86c8bb,
		24'h83e6c9,
		24'h79ddbd,
		24'h48a48e,
		24'h308479,
		24'h4eab9b,
		24'h8bf6d8,
		24'h82eac8,
		24'h7ccfb2,
		24'h98b4ab,
		24'hbc98ac,
		24'h864e72,
		24'h88699a,
		24'h612a74,
		24'h700572,
		24'h7d0078,
		24'h7d027d,
		24'h7c027e,
		24'h7c027e,
		24'h7d017e,
		24'h7f007e,
		24'h7f007e,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e017d,
		24'h7b017a,
		24'h7c007b,
		24'h820083,
		24'h840086,
		24'h7c007e,
		24'h730573,
		24'h6a1464,
		24'h2a0322,
		24'h496c45,
		24'h469544,
		24'h358138,
		24'h388043,
		24'h378e4e,
		24'h31924d,
		24'h399a4c,
		24'h399344,
		24'h479956,
		24'h236c3b,
		24'h00270c,
		24'h2e5c51,
		24'h428b85,
		24'h429490,
		24'h135b5b,
		24'h759a9d,
		24'hffffff,
		24'hbe85a4,
		24'h6d1739,
		24'h703f57,
		24'h829496,
		24'h91e3cf,
		24'h6fd6b9,
		24'h62c5ab,
		24'h27826f,
		24'h449a8e,
		24'h71cdba,
		24'h89efcf,
		24'h81e6c1,
		24'h80d8b6,
		24'h9dc8b9,
		24'h72616f,
		24'h6c406e,
		24'h4d1365,
		24'h630c76,
		24'h7b0379,
		24'h80007a,
		24'h7b037d,
		24'h7a037d,
		24'h7c027d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e017d,
		24'h7b017a,
		24'h7c007b,
		24'h820083,
		24'h840086,
		24'h7b007e,
		24'h740573,
		24'h6a1365,
		24'h2c0224,
		24'h466947,
		24'h47984d,
		24'h23702c,
		24'h3f8a4e,
		24'h368d4f,
		24'h36954f,
		24'h3c9748,
		24'h4fa151,
		24'h5ead65,
		24'h539e63,
		24'h0a3613,
		24'h305a4a,
		24'h499588,
		24'h339386,
		24'h389287,
		24'h498a86,
		24'hacc6c8,
		24'hc4bdc7,
		24'h6b656e,
		24'h5f7374,
		24'h7db9ac,
		24'h7bdcc3,
		24'h76e3c5,
		24'h72dabf,
		24'h5cbaa6,
		24'h7dd1c5,
		24'h96edd9,
		24'h8ae6c8,
		24'h86e7c2,
		24'h78dab4,
		24'h80cab2,
		24'h769697,
		24'h4e3f69,
		24'h672883,
		24'h6a0579,
		24'h80037d,
		24'h7f0079,
		24'h7b037c,
		24'h7a037c,
		24'h7c027d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007e,
		24'h7c017b,
		24'h7d007d,
		24'h820083,
		24'h840084,
		24'h7c007d,
		24'h770575,
		24'h700f6b,
		24'h30002d,
		24'h526b59,
		24'h4e9a5d,
		24'h257537,
		24'h37854a,
		24'h3c8f51,
		24'h419653,
		24'h53a057,
		24'h72b970,
		24'h76c37a,
		24'h77c485,
		24'h5d926b,
		24'h355c47,
		24'h337f6b,
		24'h42b19b,
		24'h63d1bb,
		24'h4aa794,
		24'h4d9386,
		24'h88c0b4,
		24'h6db2a2,
		24'h6fc7b0,
		24'h8bf0d4,
		24'h77e2c4,
		24'h86f3d5,
		24'h7ae5c9,
		24'h63c4af,
		24'h6dc3b4,
		24'h74c8b4,
		24'h8de3c5,
		24'h8cebc6,
		24'h7de9c1,
		24'h79e0bf,
		24'h7bc6bb,
		24'h344364,
		24'h652782,
		24'h71057a,
		24'h7f027b,
		24'h7c0076,
		24'h7c027b,
		24'h7b037b,
		24'h7c027d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h80007f,
		24'h810180,
		24'h810180,
		24'h80007f,
		24'h80007f,
		24'h80007f,
		24'h800080,
		24'h7f017e,
		24'h7f007f,
		24'h830083,
		24'h830083,
		24'h7f007f,
		24'h7a0379,
		24'h760a73,
		24'h4b0a4a,
		24'h3d4346,
		24'h48835a,
		24'h226e3a,
		24'h34844b,
		24'h3e9151,
		24'h53a360,
		24'h7ac07b,
		24'h80c47d,
		24'h76c279,
		24'h76c580,
		24'hace6b8,
		24'h406045,
		24'h11533c,
		24'h58c6ac,
		24'h65d9bd,
		24'h69d7ba,
		24'h5dbfa4,
		24'h45a188,
		24'h59c4a6,
		24'h76efcd,
		24'h84f7d7,
		24'h8bf1d5,
		24'h79dcc1,
		24'h4fb198,
		24'h2f927c,
		24'h2a8d79,
		24'h4eab94,
		24'h93eacb,
		24'h8feec9,
		24'h7febc3,
		24'h82f0cd,
		24'h75cdbf,
		24'h3e5273,
		24'h530e6a,
		24'h79057d,
		24'h7e007a,
		24'h80007a,
		24'h7d027b,
		24'h7b037b,
		24'h7d027d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h80007f,
		24'h800080,
		24'h830083,
		24'h830083,
		24'h820182,
		24'h7f017e,
		24'h7c047a,
		24'h6d156d,
		24'h14001d,
		24'h456857,
		24'h397b54,
		24'h2b7d45,
		24'h378949,
		24'h63b36e,
		24'h7dc581,
		24'h7bc17b,
		24'h7ece82,
		24'h8cde94,
		24'ha7e5b0,
		24'h345738,
		24'h18543b,
		24'h5cbba2,
		24'h66d3b5,
		24'h65d8b4,
		24'h6ad8b7,
		24'h67d1b4,
		24'h5dd6b4,
		24'h66ebc5,
		24'h81f7d6,
		24'h7edec5,
		24'h51a891,
		24'h348d76,
		24'h369983,
		24'h33a38b,
		24'h69d2b6,
		24'h8fedcb,
		24'h88e9c4,
		24'h81e9c2,
		24'h77dfbf,
		24'h4fa397,
		24'h536185,
		24'h5e0d6e,
		24'h7d027c,
		24'h7f017b,
		24'h80007b,
		24'h7f017b,
		24'h7d027b,
		24'h7e017d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810181,
		24'h810181,
		24'h820181,
		24'h820082,
		24'h820082,
		24'h820082,
		24'h820082,
		24'h820182,
		24'h820181,
		24'h740a75,
		24'h390c40,
		24'h354045,
		24'h538a6e,
		24'h20713d,
		24'h2a7e3d,
		24'h5db069,
		24'h75c37f,
		24'h73c17a,
		24'h86db8a,
		24'h94e898,
		24'h9bdda3,
		24'h64926e,
		24'h2d5c44,
		24'h5a9a85,
		24'h74cbb0,
		24'h6fd9b5,
		24'h72debc,
		24'h73dec0,
		24'h65ddbc,
		24'h5bdeb9,
		24'h7af2d0,
		24'h63caad,
		24'h2e8c73,
		24'h37937b,
		24'h40a38c,
		24'h65d0b9,
		24'h8cf1d6,
		24'h90efcc,
		24'h8ef1ca,
		24'h7ce7be,
		24'h56bd9c,
		24'h47968b,
		24'h666d92,
		24'h64096e,
		24'h81007d,
		24'h7f007c,
		24'h7f007c,
		24'h7f007c,
		24'h7f017c,
		24'h7e017d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h820082,
		24'h820082,
		24'h820082,
		24'h820082,
		24'h820082,
		24'h820082,
		24'h820082,
		24'h830083,
		24'h860086,
		24'h7b037c,
		24'h651c67,
		24'h1a0724,
		24'h4f7264,
		24'h377d51,
		24'h257537,
		24'h5aae67,
		24'h6dc47e,
		24'h68c078,
		24'h80d987,
		24'h90e593,
		24'h8fd798,
		24'hb1ebc1,
		24'h3c6048,
		24'h4a6e5e,
		24'h94d6bd,
		24'h8ae6c2,
		24'h96f7d6,
		24'h6ccbaf,
		24'h50bb9d,
		24'h63d9b7,
		24'h71e3c3,
		24'h71dbbe,
		24'h59b9a0,
		24'h5cb4a0,
		24'h72c7b9,
		24'h9bede2,
		24'h87d5c6,
		24'h6bb9a0,
		24'h76ceb0,
		24'h7ae0bd,
		24'h60c0a6,
		24'h94dad5,
		24'h63608a,
		24'h680770,
		24'h83007e,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007d,
		24'h7e017d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h820081,
		24'h820081,
		24'h820081,
		24'h820081,
		24'h820081,
		24'h820081,
		24'h820082,
		24'h830083,
		24'h850085,
		24'h80017f,
		24'h750f73,
		24'h420444,
		24'h413d4f,
		24'h59806d,
		24'h347042,
		24'h5da86a,
		24'h68c17d,
		24'h63c17a,
		24'h7cd68b,
		24'h8bdd93,
		24'h90da9c,
		24'ha2e3b3,
		24'h325e3d,
		24'h4f7962,
		24'haeefd3,
		24'h80d1af,
		24'h5fb496,
		24'h287d63,
		24'h1f775c,
		24'h57b397,
		24'h57ad95,
		24'h6cb7a7,
		24'h87bebd,
		24'h8db2bf,
		24'h91aec1,
		24'h95aec3,
		24'h73889d,
		24'h2c4453,
		24'h436e75,
		24'h84c5c5,
		24'ha9ecef,
		24'ha1d0e1,
		24'h6a5b92,
		24'h690571,
		24'h82007e,
		24'h7f007d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7e017e,
		24'h7e017e,
		24'h7f007e,
		24'h7f007e,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h820082,
		24'h820082,
		24'h810081,
		24'h820180,
		24'h7f007a,
		24'h760e73,
		24'h3a073f,
		24'h45434f,
		24'h3b5a43,
		24'h599363,
		24'h66b778,
		24'h62c07b,
		24'h79d18a,
		24'h92df9e,
		24'h7ec88c,
		24'h74bd86,
		24'h316e3f,
		24'h326941,
		24'h67a884,
		24'h4a9472,
		24'h287353,
		24'h38856a,
		24'h4a9177,
		24'h548f7a,
		24'h5b867d,
		24'h485d67,
		24'h484163,
		24'h56336b,
		24'h5e3271,
		24'h633577,
		24'h5f2f71,
		24'h4f2363,
		24'h3c2861,
		24'h444f7d,
		24'h90a6d0,
		24'h808bbb,
		24'h64408b,
		24'h6d0576,
		24'h80007e,
		24'h7e017d,
		24'h7e017d,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h820081,
		24'h820081,
		24'h810180,
		24'h810080,
		24'h880389,
		24'h7e0782,
		24'h681b6c,
		24'h1f0024,
		24'h303c35,
		24'h4b7852,
		24'h68ac73,
		24'h71c17e,
		24'h64b46b,
		24'h73be76,
		24'h68b36c,
		24'h57a25f,
		24'h5da96c,
		24'h3b7a42,
		24'h225e2b,
		24'h6ab283,
		24'ha4eebd,
		24'h9ee5b8,
		24'ha6ddbd,
		24'habcbbf,
		24'h8b8b9a,
		24'h603c68,
		24'h57185d,
		24'h5d0961,
		24'h650a6a,
		24'h670b6d,
		24'h6b0f70,
		24'h691071,
		24'h5f1974,
		24'h4a1f70,
		24'h3d1c69,
		24'h401667,
		24'h571171,
		24'h76067c,
		24'h80007e,
		24'h7e017e,
		24'h7e017e,
		24'h7f007e,
		24'h7f007e,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h810180,
		24'h800083,
		24'h80028b,
		24'h770282,
		24'h6b0f70,
		24'h2e0030,
		24'h444248,
		24'h4b6f52,
		24'h72aa75,
		24'h7cbc7a,
		24'h61a458,
		24'h4c9040,
		24'h81c679,
		24'ha3e79f,
		24'ha0e4a0,
		24'ha2e6a8,
		24'ha2e5ac,
		24'ha0e1aa,
		24'h9edea3,
		24'h99d099,
		24'h9dc0a1,
		24'h888b90,
		24'h5c2f5d,
		24'h63095b,
		24'h7c0d74,
		24'h810d7e,
		24'h800b81,
		24'h7c097d,
		24'h790679,
		24'h7a057b,
		24'h720678,
		24'h6c0d7b,
		24'h620975,
		24'h721283,
		24'h790d81,
		24'h7b017e,
		24'h80007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h800180,
		24'h7f0180,
		24'h82068a,
		24'h75007c,
		24'h751176,
		24'h40013e,
		24'h635667,
		24'h48644d,
		24'h609461,
		24'h558f4d,
		24'h77aa6d,
		24'h7fa774,
		24'h6f9566,
		24'h83aa7e,
		24'h8aaf8a,
		24'h8bae90,
		24'h93b79c,
		24'h97baa3,
		24'h9db9a2,
		24'h7c8779,
		24'h625061,
		24'h653267,
		24'h630e64,
		24'h780676,
		24'h840580,
		24'h860583,
		24'h830484,
		24'h7a017e,
		24'h77017c,
		24'h7e0281,
		24'h79007d,
		24'h7b0180,
		24'h78017e,
		24'h810684,
		24'h79007b,
		24'h7f0080,
		24'h7f0080,
		24'h7f0080,
		24'h7f0080,
		24'h7f0080,
		24'h7f0080,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7d027c,
		24'h780375,
		24'h73086b,
		24'h580851,
		24'h5d3d5e,
		24'h36463d,
		24'h507d52,
		24'h50824c,
		24'h738c6f,
		24'h5b5c59,
		24'h40393f,
		24'h423c44,
		24'h3f3846,
		24'h50485c,
		24'h655c75,
		24'h695d7c,
		24'h6d507b,
		24'h622c6a,
		24'h5c0960,
		24'h730773,
		24'h7b0782,
		24'h790284,
		24'h7d0083,
		24'h7f0082,
		24'h7e0083,
		24'h7c0185,
		24'h7b0286,
		24'h790284,
		24'h7b0082,
		24'h820083,
		24'h810084,
		24'h7f0081,
		24'h7f0082,
		24'h7f0081,
		24'h7f0081,
		24'h7f0081,
		24'h7f0081,
		24'h7e0081,
		24'h7e0081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e017e,
		24'h7d027a,
		24'h7a0478,
		24'h780776,
		24'h6e0d6c,
		24'h410041,
		24'h1c001d,
		24'h6f6a6d,
		24'h5b6055,
		24'h4d3748,
		24'h52224e,
		24'h551f52,
		24'h501a51,
		24'h511a57,
		24'h50195b,
		24'h4a1259,
		24'h541564,
		24'h62116e,
		24'h6b0571,
		24'h770379,
		24'h800380,
		24'h800284,
		24'h7e0185,
		24'h7f0086,
		24'h830086,
		24'h830085,
		24'h800084,
		24'h7c0184,
		24'h790383,
		24'h7d0082,
		24'h850082,
		24'h830082,
		24'h7d0081,
		24'h7d0081,
		24'h7f0081,
		24'h7f0081,
		24'h7f0081,
		24'h7f0081,
		24'h7e0081,
		24'h7e0081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7c027e,
		24'h7b037e,
		24'h790381,
		24'h780381,
		24'h710070,
		24'h710969,
		24'h6b2062,
		24'h602356,
		24'h621356,
		24'h700f65,
		24'h79136f,
		24'h710b6a,
		24'h730d72,
		24'h710974,
		24'h68006f,
		24'h710479,
		24'h7e0381,
		24'h850085,
		24'h7f017e,
		24'h750173,
		24'h790177,
		24'h7f007d,
		24'h840083,
		24'h850088,
		24'h870086,
		24'h860080,
		24'h81017e,
		24'h7a027e,
		24'h7e017e,
		24'h85007e,
		24'h82007e,
		24'h79037e,
		24'h79027f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7c017f,
		24'h7b0280,
		24'h7c0184,
		24'h7e0086,
		24'h80007e,
		24'h810077,
		24'h74036b,
		24'h730e6b,
		24'h76076c,
		24'h7d0472,
		24'h7e0275,
		24'h7a0074,
		24'h7c0078,
		24'h7e017d,
		24'h800283,
		24'h850689,
		24'h8a038a,
		24'h8b0088,
		24'h80007f,
		24'h7c047b,
		24'h81057e,
		24'h80007c,
		24'h830081,
		24'h840085,
		24'h860084,
		24'h86007f,
		24'h81017d,
		24'h7c027d,
		24'h7e017d,
		24'h83007d,
		24'h80017d,
		24'h79047d,
		24'h79037f,
		24'h7d017f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7c017f,
		24'h7c017f,
		24'h7e0080,
		24'h7f0080,
		24'h810080,
		24'h80007d,
		24'h7d027b,
		24'h7b0378,
		24'h7c027a,
		24'h7d007c,
		24'h7e017c,
		24'h7f017d,
		24'h7e017e,
		24'h7e007e,
		24'h7e007f,
		24'h7e007f,
		24'h800080,
		24'h820181,
		24'h800180,
		24'h7e007e,
		24'h7e007d,
		24'h80007e,
		24'h800080,
		24'h800080,
		24'h81007f,
		24'h82007f,
		24'h80007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7d017f,
		24'h7d017f,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f0080,
		24'h7f0080,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e0081,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7c017f,
		24'h7c017f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7c017f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7e007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007d,
		24'h7f007d,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007d,
		24'h81007d,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h7f007f,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007d,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h81007f,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		24'h810081,
		0x810081
	};

    always_ff @(posedge clk) begin
        o_rd_data[0][2] <= bulbasaur_rom_buf[i_rd_addr][3*bpp_p-1-:8];
        o_rd_data[0][1] <= bulbasaur_rom_buf[i_rd_addr][2*bpp_p-1-:8];
        o_rd_data[0][0] <= bulbasaur_rom_buf[i_rd_addr][1*bpp_p-1-:8];

        o_rd_data[1][2] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][3*bpp_p-1-:8];
        o_rd_data[1][1] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][2*bpp_p-1-:8];
        o_rd_data[1][0] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][1*bpp_p-1-:8];
    end
endmodule