module test_bars_rom_new #(
    parameter hpixel_p = 64,
    parameter vpixel_p = 64,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

    // Clock and reset
    input logic clk,
    input logic rst_n,

    /* Pixel read interface */
    input logic [addr_width_p-1:0] i_rd_addr,
    output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
    );


    always_ff @(posedge clk) begin
        case (i_rd_addr)
		12'd0000: rd_data_0 <= 24'hffffff;
		12'd0001: rd_data_0 <= 24'hffffff;
		12'd0002: rd_data_0 <= 24'hffffff;
		12'd0003: rd_data_0 <= 24'hffffff;
		12'd0004: rd_data_0 <= 24'hffffff;
		12'd0005: rd_data_0 <= 24'hffffff;
		12'd0006: rd_data_0 <= 24'hffffff;
		12'd0007: rd_data_0 <= 24'hffffff;
		12'd0008: rd_data_0 <= 24'hffff00;
		12'd0009: rd_data_0 <= 24'hffff00;
		12'd0010: rd_data_0 <= 24'hffff00;
		12'd0011: rd_data_0 <= 24'hffff00;
		12'd0012: rd_data_0 <= 24'hffff00;
		12'd0013: rd_data_0 <= 24'hffff00;
		12'd0014: rd_data_0 <= 24'hffff00;
		12'd0015: rd_data_0 <= 24'hffff00;
		12'd0016: rd_data_0 <= 24'h00ffff;
		12'd0017: rd_data_0 <= 24'h00ffff;
		12'd0018: rd_data_0 <= 24'h00ffff;
		12'd0019: rd_data_0 <= 24'h00ffff;
		12'd0020: rd_data_0 <= 24'h00ffff;
		12'd0021: rd_data_0 <= 24'h00ffff;
		12'd0022: rd_data_0 <= 24'h00ffff;
		12'd0023: rd_data_0 <= 24'h00ffff;
		12'd0024: rd_data_0 <= 24'h00ff00;
		12'd0025: rd_data_0 <= 24'h00ff00;
		12'd0026: rd_data_0 <= 24'h00ff00;
		12'd0027: rd_data_0 <= 24'h00ff00;
		12'd0028: rd_data_0 <= 24'h00ff00;
		12'd0029: rd_data_0 <= 24'h00ff00;
		12'd0030: rd_data_0 <= 24'h00ff00;
		12'd0031: rd_data_0 <= 24'h00ff00;
		12'd0032: rd_data_0 <= 24'hff00ff;
		12'd0033: rd_data_0 <= 24'hff00ff;
		12'd0034: rd_data_0 <= 24'hff00ff;
		12'd0035: rd_data_0 <= 24'hff00ff;
		12'd0036: rd_data_0 <= 24'hff00ff;
		12'd0037: rd_data_0 <= 24'hff00ff;
		12'd0038: rd_data_0 <= 24'hff00ff;
		12'd0039: rd_data_0 <= 24'hff00ff;
		12'd0040: rd_data_0 <= 24'hff0000;
		12'd0041: rd_data_0 <= 24'hff0000;
		12'd0042: rd_data_0 <= 24'hff0000;
		12'd0043: rd_data_0 <= 24'hff0000;
		12'd0044: rd_data_0 <= 24'hff0000;
		12'd0045: rd_data_0 <= 24'hff0000;
		12'd0046: rd_data_0 <= 24'hff0000;
		12'd0047: rd_data_0 <= 24'hff0000;
		12'd0048: rd_data_0 <= 24'h0000ff;
		12'd0049: rd_data_0 <= 24'h0000ff;
		12'd0050: rd_data_0 <= 24'h0000ff;
		12'd0051: rd_data_0 <= 24'h0000ff;
		12'd0052: rd_data_0 <= 24'h0000ff;
		12'd0053: rd_data_0 <= 24'h0000ff;
		12'd0054: rd_data_0 <= 24'h0000ff;
		12'd0055: rd_data_0 <= 24'h0000ff;
		12'd0056: rd_data_0 <= 24'h000000;
		12'd0057: rd_data_0 <= 24'h000000;
		12'd0058: rd_data_0 <= 24'h000000;
		12'd0059: rd_data_0 <= 24'h000000;
		12'd0060: rd_data_0 <= 24'h000000;
		12'd0061: rd_data_0 <= 24'h000000;
		12'd0062: rd_data_0 <= 24'h000000;
		12'd0063: rd_data_0 <= 24'h000000;
		12'd0064: rd_data_0 <= 24'hffffff;
		12'd0065: rd_data_0 <= 24'hffffff;
		12'd0066: rd_data_0 <= 24'hffffff;
		12'd0067: rd_data_0 <= 24'hffffff;
		12'd0068: rd_data_0 <= 24'hffffff;
		12'd0069: rd_data_0 <= 24'hffffff;
		12'd0070: rd_data_0 <= 24'hffffff;
		12'd0071: rd_data_0 <= 24'hffffff;
		12'd0072: rd_data_0 <= 24'hffff00;
		12'd0073: rd_data_0 <= 24'hffff00;
		12'd0074: rd_data_0 <= 24'hffff00;
		12'd0075: rd_data_0 <= 24'hffff00;
		12'd0076: rd_data_0 <= 24'hffff00;
		12'd0077: rd_data_0 <= 24'hffff00;
		12'd0078: rd_data_0 <= 24'hffff00;
		12'd0079: rd_data_0 <= 24'hffff00;
		12'd0080: rd_data_0 <= 24'h00ffff;
		12'd0081: rd_data_0 <= 24'h00ffff;
		12'd0082: rd_data_0 <= 24'h00ffff;
		12'd0083: rd_data_0 <= 24'h00ffff;
		12'd0084: rd_data_0 <= 24'h00ffff;
		12'd0085: rd_data_0 <= 24'h00ffff;
		12'd0086: rd_data_0 <= 24'h00ffff;
		12'd0087: rd_data_0 <= 24'h00ffff;
		12'd0088: rd_data_0 <= 24'h00ff00;
		12'd0089: rd_data_0 <= 24'h00ff00;
		12'd0090: rd_data_0 <= 24'h00ff00;
		12'd0091: rd_data_0 <= 24'h00ff00;
		12'd0092: rd_data_0 <= 24'h00ff00;
		12'd0093: rd_data_0 <= 24'h00ff00;
		12'd0094: rd_data_0 <= 24'h00ff00;
		12'd0095: rd_data_0 <= 24'h00ff00;
		12'd0096: rd_data_0 <= 24'hff00ff;
		12'd0097: rd_data_0 <= 24'hff00ff;
		12'd0098: rd_data_0 <= 24'hff00ff;
		12'd0099: rd_data_0 <= 24'hff00ff;
		12'd0100: rd_data_0 <= 24'hff00ff;
		12'd0101: rd_data_0 <= 24'hff00ff;
		12'd0102: rd_data_0 <= 24'hff00ff;
		12'd0103: rd_data_0 <= 24'hff00ff;
		12'd0104: rd_data_0 <= 24'hff0000;
		12'd0105: rd_data_0 <= 24'hff0000;
		12'd0106: rd_data_0 <= 24'hff0000;
		12'd0107: rd_data_0 <= 24'hff0000;
		12'd0108: rd_data_0 <= 24'hff0000;
		12'd0109: rd_data_0 <= 24'hff0000;
		12'd0110: rd_data_0 <= 24'hff0000;
		12'd0111: rd_data_0 <= 24'hff0000;
		12'd0112: rd_data_0 <= 24'h0000ff;
		12'd0113: rd_data_0 <= 24'h0000ff;
		12'd0114: rd_data_0 <= 24'h0000ff;
		12'd0115: rd_data_0 <= 24'h0000ff;
		12'd0116: rd_data_0 <= 24'h0000ff;
		12'd0117: rd_data_0 <= 24'h0000ff;
		12'd0118: rd_data_0 <= 24'h0000ff;
		12'd0119: rd_data_0 <= 24'h0000ff;
		12'd0120: rd_data_0 <= 24'h000000;
		12'd0121: rd_data_0 <= 24'h000000;
		12'd0122: rd_data_0 <= 24'h000000;
		12'd0123: rd_data_0 <= 24'h000000;
		12'd0124: rd_data_0 <= 24'h000000;
		12'd0125: rd_data_0 <= 24'h000000;
		12'd0126: rd_data_0 <= 24'h000000;
		12'd0127: rd_data_0 <= 24'h000000;
		12'd0128: rd_data_0 <= 24'hffffff;
		12'd0129: rd_data_0 <= 24'hffffff;
		12'd0130: rd_data_0 <= 24'hffffff;
		12'd0131: rd_data_0 <= 24'hffffff;
		12'd0132: rd_data_0 <= 24'hffffff;
		12'd0133: rd_data_0 <= 24'hffffff;
		12'd0134: rd_data_0 <= 24'hffffff;
		12'd0135: rd_data_0 <= 24'hffffff;
		12'd0136: rd_data_0 <= 24'hffff00;
		12'd0137: rd_data_0 <= 24'hffff00;
		12'd0138: rd_data_0 <= 24'hffff00;
		12'd0139: rd_data_0 <= 24'hffff00;
		12'd0140: rd_data_0 <= 24'hffff00;
		12'd0141: rd_data_0 <= 24'hffff00;
		12'd0142: rd_data_0 <= 24'hffff00;
		12'd0143: rd_data_0 <= 24'hffff00;
		12'd0144: rd_data_0 <= 24'h00ffff;
		12'd0145: rd_data_0 <= 24'h00ffff;
		12'd0146: rd_data_0 <= 24'h00ffff;
		12'd0147: rd_data_0 <= 24'h00ffff;
		12'd0148: rd_data_0 <= 24'h00ffff;
		12'd0149: rd_data_0 <= 24'h00ffff;
		12'd0150: rd_data_0 <= 24'h00ffff;
		12'd0151: rd_data_0 <= 24'h00ffff;
		12'd0152: rd_data_0 <= 24'h00ff00;
		12'd0153: rd_data_0 <= 24'h00ff00;
		12'd0154: rd_data_0 <= 24'h00ff00;
		12'd0155: rd_data_0 <= 24'h00ff00;
		12'd0156: rd_data_0 <= 24'h00ff00;
		12'd0157: rd_data_0 <= 24'h00ff00;
		12'd0158: rd_data_0 <= 24'h00ff00;
		12'd0159: rd_data_0 <= 24'h00ff00;
		12'd0160: rd_data_0 <= 24'hff00ff;
		12'd0161: rd_data_0 <= 24'hff00ff;
		12'd0162: rd_data_0 <= 24'hff00ff;
		12'd0163: rd_data_0 <= 24'hff00ff;
		12'd0164: rd_data_0 <= 24'hff00ff;
		12'd0165: rd_data_0 <= 24'hff00ff;
		12'd0166: rd_data_0 <= 24'hff00ff;
		12'd0167: rd_data_0 <= 24'hff00ff;
		12'd0168: rd_data_0 <= 24'hff0000;
		12'd0169: rd_data_0 <= 24'hff0000;
		12'd0170: rd_data_0 <= 24'hff0000;
		12'd0171: rd_data_0 <= 24'hff0000;
		12'd0172: rd_data_0 <= 24'hff0000;
		12'd0173: rd_data_0 <= 24'hff0000;
		12'd0174: rd_data_0 <= 24'hff0000;
		12'd0175: rd_data_0 <= 24'hff0000;
		12'd0176: rd_data_0 <= 24'h0000ff;
		12'd0177: rd_data_0 <= 24'h0000ff;
		12'd0178: rd_data_0 <= 24'h0000ff;
		12'd0179: rd_data_0 <= 24'h0000ff;
		12'd0180: rd_data_0 <= 24'h0000ff;
		12'd0181: rd_data_0 <= 24'h0000ff;
		12'd0182: rd_data_0 <= 24'h0000ff;
		12'd0183: rd_data_0 <= 24'h0000ff;
		12'd0184: rd_data_0 <= 24'h000000;
		12'd0185: rd_data_0 <= 24'h000000;
		12'd0186: rd_data_0 <= 24'h000000;
		12'd0187: rd_data_0 <= 24'h000000;
		12'd0188: rd_data_0 <= 24'h000000;
		12'd0189: rd_data_0 <= 24'h000000;
		12'd0190: rd_data_0 <= 24'h000000;
		12'd0191: rd_data_0 <= 24'h000000;
		12'd0192: rd_data_0 <= 24'hffffff;
		12'd0193: rd_data_0 <= 24'hffffff;
		12'd0194: rd_data_0 <= 24'hffffff;
		12'd0195: rd_data_0 <= 24'hffffff;
		12'd0196: rd_data_0 <= 24'hffffff;
		12'd0197: rd_data_0 <= 24'hffffff;
		12'd0198: rd_data_0 <= 24'hffffff;
		12'd0199: rd_data_0 <= 24'hffffff;
		12'd0200: rd_data_0 <= 24'hffff00;
		12'd0201: rd_data_0 <= 24'hffff00;
		12'd0202: rd_data_0 <= 24'hffff00;
		12'd0203: rd_data_0 <= 24'hffff00;
		12'd0204: rd_data_0 <= 24'hffff00;
		12'd0205: rd_data_0 <= 24'hffff00;
		12'd0206: rd_data_0 <= 24'hffff00;
		12'd0207: rd_data_0 <= 24'hffff00;
		12'd0208: rd_data_0 <= 24'h00ffff;
		12'd0209: rd_data_0 <= 24'h00ffff;
		12'd0210: rd_data_0 <= 24'h00ffff;
		12'd0211: rd_data_0 <= 24'h00ffff;
		12'd0212: rd_data_0 <= 24'h00ffff;
		12'd0213: rd_data_0 <= 24'h00ffff;
		12'd0214: rd_data_0 <= 24'h00ffff;
		12'd0215: rd_data_0 <= 24'h00ffff;
		12'd0216: rd_data_0 <= 24'h00ff00;
		12'd0217: rd_data_0 <= 24'h00ff00;
		12'd0218: rd_data_0 <= 24'h00ff00;
		12'd0219: rd_data_0 <= 24'h00ff00;
		12'd0220: rd_data_0 <= 24'h00ff00;
		12'd0221: rd_data_0 <= 24'h00ff00;
		12'd0222: rd_data_0 <= 24'h00ff00;
		12'd0223: rd_data_0 <= 24'h00ff00;
		12'd0224: rd_data_0 <= 24'hff00ff;
		12'd0225: rd_data_0 <= 24'hff00ff;
		12'd0226: rd_data_0 <= 24'hff00ff;
		12'd0227: rd_data_0 <= 24'hff00ff;
		12'd0228: rd_data_0 <= 24'hff00ff;
		12'd0229: rd_data_0 <= 24'hff00ff;
		12'd0230: rd_data_0 <= 24'hff00ff;
		12'd0231: rd_data_0 <= 24'hff00ff;
		12'd0232: rd_data_0 <= 24'hff0000;
		12'd0233: rd_data_0 <= 24'hff0000;
		12'd0234: rd_data_0 <= 24'hff0000;
		12'd0235: rd_data_0 <= 24'hff0000;
		12'd0236: rd_data_0 <= 24'hff0000;
		12'd0237: rd_data_0 <= 24'hff0000;
		12'd0238: rd_data_0 <= 24'hff0000;
		12'd0239: rd_data_0 <= 24'hff0000;
		12'd0240: rd_data_0 <= 24'h0000ff;
		12'd0241: rd_data_0 <= 24'h0000ff;
		12'd0242: rd_data_0 <= 24'h0000ff;
		12'd0243: rd_data_0 <= 24'h0000ff;
		12'd0244: rd_data_0 <= 24'h0000ff;
		12'd0245: rd_data_0 <= 24'h0000ff;
		12'd0246: rd_data_0 <= 24'h0000ff;
		12'd0247: rd_data_0 <= 24'h0000ff;
		12'd0248: rd_data_0 <= 24'h000000;
		12'd0249: rd_data_0 <= 24'h000000;
		12'd0250: rd_data_0 <= 24'h000000;
		12'd0251: rd_data_0 <= 24'h000000;
		12'd0252: rd_data_0 <= 24'h000000;
		12'd0253: rd_data_0 <= 24'h000000;
		12'd0254: rd_data_0 <= 24'h000000;
		12'd0255: rd_data_0 <= 24'h000000;
		12'd0256: rd_data_0 <= 24'hffffff;
		12'd0257: rd_data_0 <= 24'hffffff;
		12'd0258: rd_data_0 <= 24'hffffff;
		12'd0259: rd_data_0 <= 24'hffffff;
		12'd0260: rd_data_0 <= 24'hffffff;
		12'd0261: rd_data_0 <= 24'hffffff;
		12'd0262: rd_data_0 <= 24'hffffff;
		12'd0263: rd_data_0 <= 24'hffffff;
		12'd0264: rd_data_0 <= 24'hffff00;
		12'd0265: rd_data_0 <= 24'hffff00;
		12'd0266: rd_data_0 <= 24'hffff00;
		12'd0267: rd_data_0 <= 24'hffff00;
		12'd0268: rd_data_0 <= 24'hffff00;
		12'd0269: rd_data_0 <= 24'hffff00;
		12'd0270: rd_data_0 <= 24'hffff00;
		12'd0271: rd_data_0 <= 24'hffff00;
		12'd0272: rd_data_0 <= 24'h00ffff;
		12'd0273: rd_data_0 <= 24'h00ffff;
		12'd0274: rd_data_0 <= 24'h00ffff;
		12'd0275: rd_data_0 <= 24'h00ffff;
		12'd0276: rd_data_0 <= 24'h00ffff;
		12'd0277: rd_data_0 <= 24'h00ffff;
		12'd0278: rd_data_0 <= 24'h00ffff;
		12'd0279: rd_data_0 <= 24'h00ffff;
		12'd0280: rd_data_0 <= 24'h00ff00;
		12'd0281: rd_data_0 <= 24'h00ff00;
		12'd0282: rd_data_0 <= 24'h00ff00;
		12'd0283: rd_data_0 <= 24'h00ff00;
		12'd0284: rd_data_0 <= 24'h00ff00;
		12'd0285: rd_data_0 <= 24'h00ff00;
		12'd0286: rd_data_0 <= 24'h00ff00;
		12'd0287: rd_data_0 <= 24'h00ff00;
		12'd0288: rd_data_0 <= 24'hff00ff;
		12'd0289: rd_data_0 <= 24'hff00ff;
		12'd0290: rd_data_0 <= 24'hff00ff;
		12'd0291: rd_data_0 <= 24'hff00ff;
		12'd0292: rd_data_0 <= 24'hff00ff;
		12'd0293: rd_data_0 <= 24'hff00ff;
		12'd0294: rd_data_0 <= 24'hff00ff;
		12'd0295: rd_data_0 <= 24'hff00ff;
		12'd0296: rd_data_0 <= 24'hff0000;
		12'd0297: rd_data_0 <= 24'hff0000;
		12'd0298: rd_data_0 <= 24'hff0000;
		12'd0299: rd_data_0 <= 24'hff0000;
		12'd0300: rd_data_0 <= 24'hff0000;
		12'd0301: rd_data_0 <= 24'hff0000;
		12'd0302: rd_data_0 <= 24'hff0000;
		12'd0303: rd_data_0 <= 24'hff0000;
		12'd0304: rd_data_0 <= 24'h0000ff;
		12'd0305: rd_data_0 <= 24'h0000ff;
		12'd0306: rd_data_0 <= 24'h0000ff;
		12'd0307: rd_data_0 <= 24'h0000ff;
		12'd0308: rd_data_0 <= 24'h0000ff;
		12'd0309: rd_data_0 <= 24'h0000ff;
		12'd0310: rd_data_0 <= 24'h0000ff;
		12'd0311: rd_data_0 <= 24'h0000ff;
		12'd0312: rd_data_0 <= 24'h000000;
		12'd0313: rd_data_0 <= 24'h000000;
		12'd0314: rd_data_0 <= 24'h000000;
		12'd0315: rd_data_0 <= 24'h000000;
		12'd0316: rd_data_0 <= 24'h000000;
		12'd0317: rd_data_0 <= 24'h000000;
		12'd0318: rd_data_0 <= 24'h000000;
		12'd0319: rd_data_0 <= 24'h000000;
		12'd0320: rd_data_0 <= 24'hffffff;
		12'd0321: rd_data_0 <= 24'hffffff;
		12'd0322: rd_data_0 <= 24'hffffff;
		12'd0323: rd_data_0 <= 24'hffffff;
		12'd0324: rd_data_0 <= 24'hffffff;
		12'd0325: rd_data_0 <= 24'hffffff;
		12'd0326: rd_data_0 <= 24'hffffff;
		12'd0327: rd_data_0 <= 24'hffffff;
		12'd0328: rd_data_0 <= 24'hffff00;
		12'd0329: rd_data_0 <= 24'hffff00;
		12'd0330: rd_data_0 <= 24'hffff00;
		12'd0331: rd_data_0 <= 24'hffff00;
		12'd0332: rd_data_0 <= 24'hffff00;
		12'd0333: rd_data_0 <= 24'hffff00;
		12'd0334: rd_data_0 <= 24'hffff00;
		12'd0335: rd_data_0 <= 24'hffff00;
		12'd0336: rd_data_0 <= 24'h00ffff;
		12'd0337: rd_data_0 <= 24'h00ffff;
		12'd0338: rd_data_0 <= 24'h00ffff;
		12'd0339: rd_data_0 <= 24'h00ffff;
		12'd0340: rd_data_0 <= 24'h00ffff;
		12'd0341: rd_data_0 <= 24'h00ffff;
		12'd0342: rd_data_0 <= 24'h00ffff;
		12'd0343: rd_data_0 <= 24'h00ffff;
		12'd0344: rd_data_0 <= 24'h00ff00;
		12'd0345: rd_data_0 <= 24'h00ff00;
		12'd0346: rd_data_0 <= 24'h00ff00;
		12'd0347: rd_data_0 <= 24'h00ff00;
		12'd0348: rd_data_0 <= 24'h00ff00;
		12'd0349: rd_data_0 <= 24'h00ff00;
		12'd0350: rd_data_0 <= 24'h00ff00;
		12'd0351: rd_data_0 <= 24'h00ff00;
		12'd0352: rd_data_0 <= 24'hff00ff;
		12'd0353: rd_data_0 <= 24'hff00ff;
		12'd0354: rd_data_0 <= 24'hff00ff;
		12'd0355: rd_data_0 <= 24'hff00ff;
		12'd0356: rd_data_0 <= 24'hff00ff;
		12'd0357: rd_data_0 <= 24'hff00ff;
		12'd0358: rd_data_0 <= 24'hff00ff;
		12'd0359: rd_data_0 <= 24'hff00ff;
		12'd0360: rd_data_0 <= 24'hff0000;
		12'd0361: rd_data_0 <= 24'hff0000;
		12'd0362: rd_data_0 <= 24'hff0000;
		12'd0363: rd_data_0 <= 24'hff0000;
		12'd0364: rd_data_0 <= 24'hff0000;
		12'd0365: rd_data_0 <= 24'hff0000;
		12'd0366: rd_data_0 <= 24'hff0000;
		12'd0367: rd_data_0 <= 24'hff0000;
		12'd0368: rd_data_0 <= 24'h0000ff;
		12'd0369: rd_data_0 <= 24'h0000ff;
		12'd0370: rd_data_0 <= 24'h0000ff;
		12'd0371: rd_data_0 <= 24'h0000ff;
		12'd0372: rd_data_0 <= 24'h0000ff;
		12'd0373: rd_data_0 <= 24'h0000ff;
		12'd0374: rd_data_0 <= 24'h0000ff;
		12'd0375: rd_data_0 <= 24'h0000ff;
		12'd0376: rd_data_0 <= 24'h000000;
		12'd0377: rd_data_0 <= 24'h000000;
		12'd0378: rd_data_0 <= 24'h000000;
		12'd0379: rd_data_0 <= 24'h000000;
		12'd0380: rd_data_0 <= 24'h000000;
		12'd0381: rd_data_0 <= 24'h000000;
		12'd0382: rd_data_0 <= 24'h000000;
		12'd0383: rd_data_0 <= 24'h000000;
		12'd0384: rd_data_0 <= 24'hffffff;
		12'd0385: rd_data_0 <= 24'hffffff;
		12'd0386: rd_data_0 <= 24'hffffff;
		12'd0387: rd_data_0 <= 24'hffffff;
		12'd0388: rd_data_0 <= 24'hffffff;
		12'd0389: rd_data_0 <= 24'hffffff;
		12'd0390: rd_data_0 <= 24'hffffff;
		12'd0391: rd_data_0 <= 24'hffffff;
		12'd0392: rd_data_0 <= 24'hffff00;
		12'd0393: rd_data_0 <= 24'hffff00;
		12'd0394: rd_data_0 <= 24'hffff00;
		12'd0395: rd_data_0 <= 24'hffff00;
		12'd0396: rd_data_0 <= 24'hffff00;
		12'd0397: rd_data_0 <= 24'hffff00;
		12'd0398: rd_data_0 <= 24'hffff00;
		12'd0399: rd_data_0 <= 24'hffff00;
		12'd0400: rd_data_0 <= 24'h00ffff;
		12'd0401: rd_data_0 <= 24'h00ffff;
		12'd0402: rd_data_0 <= 24'h00ffff;
		12'd0403: rd_data_0 <= 24'h00ffff;
		12'd0404: rd_data_0 <= 24'h00ffff;
		12'd0405: rd_data_0 <= 24'h00ffff;
		12'd0406: rd_data_0 <= 24'h00ffff;
		12'd0407: rd_data_0 <= 24'h00ffff;
		12'd0408: rd_data_0 <= 24'h00ff00;
		12'd0409: rd_data_0 <= 24'h00ff00;
		12'd0410: rd_data_0 <= 24'h00ff00;
		12'd0411: rd_data_0 <= 24'h00ff00;
		12'd0412: rd_data_0 <= 24'h00ff00;
		12'd0413: rd_data_0 <= 24'h00ff00;
		12'd0414: rd_data_0 <= 24'h00ff00;
		12'd0415: rd_data_0 <= 24'h00ff00;
		12'd0416: rd_data_0 <= 24'hff00ff;
		12'd0417: rd_data_0 <= 24'hff00ff;
		12'd0418: rd_data_0 <= 24'hff00ff;
		12'd0419: rd_data_0 <= 24'hff00ff;
		12'd0420: rd_data_0 <= 24'hff00ff;
		12'd0421: rd_data_0 <= 24'hff00ff;
		12'd0422: rd_data_0 <= 24'hff00ff;
		12'd0423: rd_data_0 <= 24'hff00ff;
		12'd0424: rd_data_0 <= 24'hff0000;
		12'd0425: rd_data_0 <= 24'hff0000;
		12'd0426: rd_data_0 <= 24'hff0000;
		12'd0427: rd_data_0 <= 24'hff0000;
		12'd0428: rd_data_0 <= 24'hff0000;
		12'd0429: rd_data_0 <= 24'hff0000;
		12'd0430: rd_data_0 <= 24'hff0000;
		12'd0431: rd_data_0 <= 24'hff0000;
		12'd0432: rd_data_0 <= 24'h0000ff;
		12'd0433: rd_data_0 <= 24'h0000ff;
		12'd0434: rd_data_0 <= 24'h0000ff;
		12'd0435: rd_data_0 <= 24'h0000ff;
		12'd0436: rd_data_0 <= 24'h0000ff;
		12'd0437: rd_data_0 <= 24'h0000ff;
		12'd0438: rd_data_0 <= 24'h0000ff;
		12'd0439: rd_data_0 <= 24'h0000ff;
		12'd0440: rd_data_0 <= 24'h000000;
		12'd0441: rd_data_0 <= 24'h000000;
		12'd0442: rd_data_0 <= 24'h000000;
		12'd0443: rd_data_0 <= 24'h000000;
		12'd0444: rd_data_0 <= 24'h000000;
		12'd0445: rd_data_0 <= 24'h000000;
		12'd0446: rd_data_0 <= 24'h000000;
		12'd0447: rd_data_0 <= 24'h000000;
		12'd0448: rd_data_0 <= 24'hffffff;
		12'd0449: rd_data_0 <= 24'hffffff;
		12'd0450: rd_data_0 <= 24'hffffff;
		12'd0451: rd_data_0 <= 24'hffffff;
		12'd0452: rd_data_0 <= 24'hffffff;
		12'd0453: rd_data_0 <= 24'hffffff;
		12'd0454: rd_data_0 <= 24'hffffff;
		12'd0455: rd_data_0 <= 24'hffffff;
		12'd0456: rd_data_0 <= 24'hffff00;
		12'd0457: rd_data_0 <= 24'hffff00;
		12'd0458: rd_data_0 <= 24'hffff00;
		12'd0459: rd_data_0 <= 24'hffff00;
		12'd0460: rd_data_0 <= 24'hffff00;
		12'd0461: rd_data_0 <= 24'hffff00;
		12'd0462: rd_data_0 <= 24'hffff00;
		12'd0463: rd_data_0 <= 24'hffff00;
		12'd0464: rd_data_0 <= 24'h00ffff;
		12'd0465: rd_data_0 <= 24'h00ffff;
		12'd0466: rd_data_0 <= 24'h00ffff;
		12'd0467: rd_data_0 <= 24'h00ffff;
		12'd0468: rd_data_0 <= 24'h00ffff;
		12'd0469: rd_data_0 <= 24'h00ffff;
		12'd0470: rd_data_0 <= 24'h00ffff;
		12'd0471: rd_data_0 <= 24'h00ffff;
		12'd0472: rd_data_0 <= 24'h00ff00;
		12'd0473: rd_data_0 <= 24'h00ff00;
		12'd0474: rd_data_0 <= 24'h00ff00;
		12'd0475: rd_data_0 <= 24'h00ff00;
		12'd0476: rd_data_0 <= 24'h00ff00;
		12'd0477: rd_data_0 <= 24'h00ff00;
		12'd0478: rd_data_0 <= 24'h00ff00;
		12'd0479: rd_data_0 <= 24'h00ff00;
		12'd0480: rd_data_0 <= 24'hff00ff;
		12'd0481: rd_data_0 <= 24'hff00ff;
		12'd0482: rd_data_0 <= 24'hff00ff;
		12'd0483: rd_data_0 <= 24'hff00ff;
		12'd0484: rd_data_0 <= 24'hff00ff;
		12'd0485: rd_data_0 <= 24'hff00ff;
		12'd0486: rd_data_0 <= 24'hff00ff;
		12'd0487: rd_data_0 <= 24'hff00ff;
		12'd0488: rd_data_0 <= 24'hff0000;
		12'd0489: rd_data_0 <= 24'hff0000;
		12'd0490: rd_data_0 <= 24'hff0000;
		12'd0491: rd_data_0 <= 24'hff0000;
		12'd0492: rd_data_0 <= 24'hff0000;
		12'd0493: rd_data_0 <= 24'hff0000;
		12'd0494: rd_data_0 <= 24'hff0000;
		12'd0495: rd_data_0 <= 24'hff0000;
		12'd0496: rd_data_0 <= 24'h0000ff;
		12'd0497: rd_data_0 <= 24'h0000ff;
		12'd0498: rd_data_0 <= 24'h0000ff;
		12'd0499: rd_data_0 <= 24'h0000ff;
		12'd0500: rd_data_0 <= 24'h0000ff;
		12'd0501: rd_data_0 <= 24'h0000ff;
		12'd0502: rd_data_0 <= 24'h0000ff;
		12'd0503: rd_data_0 <= 24'h0000ff;
		12'd0504: rd_data_0 <= 24'h000000;
		12'd0505: rd_data_0 <= 24'h000000;
		12'd0506: rd_data_0 <= 24'h000000;
		12'd0507: rd_data_0 <= 24'h000000;
		12'd0508: rd_data_0 <= 24'h000000;
		12'd0509: rd_data_0 <= 24'h000000;
		12'd0510: rd_data_0 <= 24'h000000;
		12'd0511: rd_data_0 <= 24'h000000;
		12'd0512: rd_data_0 <= 24'hffffff;
		12'd0513: rd_data_0 <= 24'hffffff;
		12'd0514: rd_data_0 <= 24'hffffff;
		12'd0515: rd_data_0 <= 24'hffffff;
		12'd0516: rd_data_0 <= 24'hffffff;
		12'd0517: rd_data_0 <= 24'hffffff;
		12'd0518: rd_data_0 <= 24'hffffff;
		12'd0519: rd_data_0 <= 24'hffffff;
		12'd0520: rd_data_0 <= 24'hffff00;
		12'd0521: rd_data_0 <= 24'hffff00;
		12'd0522: rd_data_0 <= 24'hffff00;
		12'd0523: rd_data_0 <= 24'hffff00;
		12'd0524: rd_data_0 <= 24'hffff00;
		12'd0525: rd_data_0 <= 24'hffff00;
		12'd0526: rd_data_0 <= 24'hffff00;
		12'd0527: rd_data_0 <= 24'hffff00;
		12'd0528: rd_data_0 <= 24'h00ffff;
		12'd0529: rd_data_0 <= 24'h00ffff;
		12'd0530: rd_data_0 <= 24'h00ffff;
		12'd0531: rd_data_0 <= 24'h00ffff;
		12'd0532: rd_data_0 <= 24'h00ffff;
		12'd0533: rd_data_0 <= 24'h00ffff;
		12'd0534: rd_data_0 <= 24'h00ffff;
		12'd0535: rd_data_0 <= 24'h00ffff;
		12'd0536: rd_data_0 <= 24'h00ff00;
		12'd0537: rd_data_0 <= 24'h00ff00;
		12'd0538: rd_data_0 <= 24'h00ff00;
		12'd0539: rd_data_0 <= 24'h00ff00;
		12'd0540: rd_data_0 <= 24'h00ff00;
		12'd0541: rd_data_0 <= 24'h00ff00;
		12'd0542: rd_data_0 <= 24'h00ff00;
		12'd0543: rd_data_0 <= 24'h00ff00;
		12'd0544: rd_data_0 <= 24'hff00ff;
		12'd0545: rd_data_0 <= 24'hff00ff;
		12'd0546: rd_data_0 <= 24'hff00ff;
		12'd0547: rd_data_0 <= 24'hff00ff;
		12'd0548: rd_data_0 <= 24'hff00ff;
		12'd0549: rd_data_0 <= 24'hff00ff;
		12'd0550: rd_data_0 <= 24'hff00ff;
		12'd0551: rd_data_0 <= 24'hff00ff;
		12'd0552: rd_data_0 <= 24'hff0000;
		12'd0553: rd_data_0 <= 24'hff0000;
		12'd0554: rd_data_0 <= 24'hff0000;
		12'd0555: rd_data_0 <= 24'hff0000;
		12'd0556: rd_data_0 <= 24'hff0000;
		12'd0557: rd_data_0 <= 24'hff0000;
		12'd0558: rd_data_0 <= 24'hff0000;
		12'd0559: rd_data_0 <= 24'hff0000;
		12'd0560: rd_data_0 <= 24'h0000ff;
		12'd0561: rd_data_0 <= 24'h0000ff;
		12'd0562: rd_data_0 <= 24'h0000ff;
		12'd0563: rd_data_0 <= 24'h0000ff;
		12'd0564: rd_data_0 <= 24'h0000ff;
		12'd0565: rd_data_0 <= 24'h0000ff;
		12'd0566: rd_data_0 <= 24'h0000ff;
		12'd0567: rd_data_0 <= 24'h0000ff;
		12'd0568: rd_data_0 <= 24'h000000;
		12'd0569: rd_data_0 <= 24'h000000;
		12'd0570: rd_data_0 <= 24'h000000;
		12'd0571: rd_data_0 <= 24'h000000;
		12'd0572: rd_data_0 <= 24'h000000;
		12'd0573: rd_data_0 <= 24'h000000;
		12'd0574: rd_data_0 <= 24'h000000;
		12'd0575: rd_data_0 <= 24'h000000;
		12'd0576: rd_data_0 <= 24'hffffff;
		12'd0577: rd_data_0 <= 24'hffffff;
		12'd0578: rd_data_0 <= 24'hffffff;
		12'd0579: rd_data_0 <= 24'hffffff;
		12'd0580: rd_data_0 <= 24'hffffff;
		12'd0581: rd_data_0 <= 24'hffffff;
		12'd0582: rd_data_0 <= 24'hffffff;
		12'd0583: rd_data_0 <= 24'hffffff;
		12'd0584: rd_data_0 <= 24'hffff00;
		12'd0585: rd_data_0 <= 24'hffff00;
		12'd0586: rd_data_0 <= 24'hffff00;
		12'd0587: rd_data_0 <= 24'hffff00;
		12'd0588: rd_data_0 <= 24'hffff00;
		12'd0589: rd_data_0 <= 24'hffff00;
		12'd0590: rd_data_0 <= 24'hffff00;
		12'd0591: rd_data_0 <= 24'hffff00;
		12'd0592: rd_data_0 <= 24'h00ffff;
		12'd0593: rd_data_0 <= 24'h00ffff;
		12'd0594: rd_data_0 <= 24'h00ffff;
		12'd0595: rd_data_0 <= 24'h00ffff;
		12'd0596: rd_data_0 <= 24'h00ffff;
		12'd0597: rd_data_0 <= 24'h00ffff;
		12'd0598: rd_data_0 <= 24'h00ffff;
		12'd0599: rd_data_0 <= 24'h00ffff;
		12'd0600: rd_data_0 <= 24'h00ff00;
		12'd0601: rd_data_0 <= 24'h00ff00;
		12'd0602: rd_data_0 <= 24'h00ff00;
		12'd0603: rd_data_0 <= 24'h00ff00;
		12'd0604: rd_data_0 <= 24'h00ff00;
		12'd0605: rd_data_0 <= 24'h00ff00;
		12'd0606: rd_data_0 <= 24'h00ff00;
		12'd0607: rd_data_0 <= 24'h00ff00;
		12'd0608: rd_data_0 <= 24'hff00ff;
		12'd0609: rd_data_0 <= 24'hff00ff;
		12'd0610: rd_data_0 <= 24'hff00ff;
		12'd0611: rd_data_0 <= 24'hff00ff;
		12'd0612: rd_data_0 <= 24'hff00ff;
		12'd0613: rd_data_0 <= 24'hff00ff;
		12'd0614: rd_data_0 <= 24'hff00ff;
		12'd0615: rd_data_0 <= 24'hff00ff;
		12'd0616: rd_data_0 <= 24'hff0000;
		12'd0617: rd_data_0 <= 24'hff0000;
		12'd0618: rd_data_0 <= 24'hff0000;
		12'd0619: rd_data_0 <= 24'hff0000;
		12'd0620: rd_data_0 <= 24'hff0000;
		12'd0621: rd_data_0 <= 24'hff0000;
		12'd0622: rd_data_0 <= 24'hff0000;
		12'd0623: rd_data_0 <= 24'hff0000;
		12'd0624: rd_data_0 <= 24'h0000ff;
		12'd0625: rd_data_0 <= 24'h0000ff;
		12'd0626: rd_data_0 <= 24'h0000ff;
		12'd0627: rd_data_0 <= 24'h0000ff;
		12'd0628: rd_data_0 <= 24'h0000ff;
		12'd0629: rd_data_0 <= 24'h0000ff;
		12'd0630: rd_data_0 <= 24'h0000ff;
		12'd0631: rd_data_0 <= 24'h0000ff;
		12'd0632: rd_data_0 <= 24'h000000;
		12'd0633: rd_data_0 <= 24'h000000;
		12'd0634: rd_data_0 <= 24'h000000;
		12'd0635: rd_data_0 <= 24'h000000;
		12'd0636: rd_data_0 <= 24'h000000;
		12'd0637: rd_data_0 <= 24'h000000;
		12'd0638: rd_data_0 <= 24'h000000;
		12'd0639: rd_data_0 <= 24'h000000;
		12'd0640: rd_data_0 <= 24'hffffff;
		12'd0641: rd_data_0 <= 24'hffffff;
		12'd0642: rd_data_0 <= 24'hffffff;
		12'd0643: rd_data_0 <= 24'hffffff;
		12'd0644: rd_data_0 <= 24'hffffff;
		12'd0645: rd_data_0 <= 24'hffffff;
		12'd0646: rd_data_0 <= 24'hffffff;
		12'd0647: rd_data_0 <= 24'hffffff;
		12'd0648: rd_data_0 <= 24'hffff00;
		12'd0649: rd_data_0 <= 24'hffff00;
		12'd0650: rd_data_0 <= 24'hffff00;
		12'd0651: rd_data_0 <= 24'hffff00;
		12'd0652: rd_data_0 <= 24'hffff00;
		12'd0653: rd_data_0 <= 24'hffff00;
		12'd0654: rd_data_0 <= 24'hffff00;
		12'd0655: rd_data_0 <= 24'hffff00;
		12'd0656: rd_data_0 <= 24'h00ffff;
		12'd0657: rd_data_0 <= 24'h00ffff;
		12'd0658: rd_data_0 <= 24'h00ffff;
		12'd0659: rd_data_0 <= 24'h00ffff;
		12'd0660: rd_data_0 <= 24'h00ffff;
		12'd0661: rd_data_0 <= 24'h00ffff;
		12'd0662: rd_data_0 <= 24'h00ffff;
		12'd0663: rd_data_0 <= 24'h00ffff;
		12'd0664: rd_data_0 <= 24'h00ff00;
		12'd0665: rd_data_0 <= 24'h00ff00;
		12'd0666: rd_data_0 <= 24'h00ff00;
		12'd0667: rd_data_0 <= 24'h00ff00;
		12'd0668: rd_data_0 <= 24'h00ff00;
		12'd0669: rd_data_0 <= 24'h00ff00;
		12'd0670: rd_data_0 <= 24'h00ff00;
		12'd0671: rd_data_0 <= 24'h00ff00;
		12'd0672: rd_data_0 <= 24'hff00ff;
		12'd0673: rd_data_0 <= 24'hff00ff;
		12'd0674: rd_data_0 <= 24'hff00ff;
		12'd0675: rd_data_0 <= 24'hff00ff;
		12'd0676: rd_data_0 <= 24'hff00ff;
		12'd0677: rd_data_0 <= 24'hff00ff;
		12'd0678: rd_data_0 <= 24'hff00ff;
		12'd0679: rd_data_0 <= 24'hff00ff;
		12'd0680: rd_data_0 <= 24'hff0000;
		12'd0681: rd_data_0 <= 24'hff0000;
		12'd0682: rd_data_0 <= 24'hff0000;
		12'd0683: rd_data_0 <= 24'hff0000;
		12'd0684: rd_data_0 <= 24'hff0000;
		12'd0685: rd_data_0 <= 24'hff0000;
		12'd0686: rd_data_0 <= 24'hff0000;
		12'd0687: rd_data_0 <= 24'hff0000;
		12'd0688: rd_data_0 <= 24'h0000ff;
		12'd0689: rd_data_0 <= 24'h0000ff;
		12'd0690: rd_data_0 <= 24'h0000ff;
		12'd0691: rd_data_0 <= 24'h0000ff;
		12'd0692: rd_data_0 <= 24'h0000ff;
		12'd0693: rd_data_0 <= 24'h0000ff;
		12'd0694: rd_data_0 <= 24'h0000ff;
		12'd0695: rd_data_0 <= 24'h0000ff;
		12'd0696: rd_data_0 <= 24'h000000;
		12'd0697: rd_data_0 <= 24'h000000;
		12'd0698: rd_data_0 <= 24'h000000;
		12'd0699: rd_data_0 <= 24'h000000;
		12'd0700: rd_data_0 <= 24'h000000;
		12'd0701: rd_data_0 <= 24'h000000;
		12'd0702: rd_data_0 <= 24'h000000;
		12'd0703: rd_data_0 <= 24'h000000;
		12'd0704: rd_data_0 <= 24'hffffff;
		12'd0705: rd_data_0 <= 24'hffffff;
		12'd0706: rd_data_0 <= 24'hffffff;
		12'd0707: rd_data_0 <= 24'hffffff;
		12'd0708: rd_data_0 <= 24'hffffff;
		12'd0709: rd_data_0 <= 24'hffffff;
		12'd0710: rd_data_0 <= 24'hffffff;
		12'd0711: rd_data_0 <= 24'hffffff;
		12'd0712: rd_data_0 <= 24'hffff00;
		12'd0713: rd_data_0 <= 24'hffff00;
		12'd0714: rd_data_0 <= 24'hffff00;
		12'd0715: rd_data_0 <= 24'hffff00;
		12'd0716: rd_data_0 <= 24'hffff00;
		12'd0717: rd_data_0 <= 24'hffff00;
		12'd0718: rd_data_0 <= 24'hffff00;
		12'd0719: rd_data_0 <= 24'hffff00;
		12'd0720: rd_data_0 <= 24'h00ffff;
		12'd0721: rd_data_0 <= 24'h00ffff;
		12'd0722: rd_data_0 <= 24'h00ffff;
		12'd0723: rd_data_0 <= 24'h00ffff;
		12'd0724: rd_data_0 <= 24'h00ffff;
		12'd0725: rd_data_0 <= 24'h00ffff;
		12'd0726: rd_data_0 <= 24'h00ffff;
		12'd0727: rd_data_0 <= 24'h00ffff;
		12'd0728: rd_data_0 <= 24'h00ff00;
		12'd0729: rd_data_0 <= 24'h00ff00;
		12'd0730: rd_data_0 <= 24'h00ff00;
		12'd0731: rd_data_0 <= 24'h00ff00;
		12'd0732: rd_data_0 <= 24'h00ff00;
		12'd0733: rd_data_0 <= 24'h00ff00;
		12'd0734: rd_data_0 <= 24'h00ff00;
		12'd0735: rd_data_0 <= 24'h00ff00;
		12'd0736: rd_data_0 <= 24'hff00ff;
		12'd0737: rd_data_0 <= 24'hff00ff;
		12'd0738: rd_data_0 <= 24'hff00ff;
		12'd0739: rd_data_0 <= 24'hff00ff;
		12'd0740: rd_data_0 <= 24'hff00ff;
		12'd0741: rd_data_0 <= 24'hff00ff;
		12'd0742: rd_data_0 <= 24'hff00ff;
		12'd0743: rd_data_0 <= 24'hff00ff;
		12'd0744: rd_data_0 <= 24'hff0000;
		12'd0745: rd_data_0 <= 24'hff0000;
		12'd0746: rd_data_0 <= 24'hff0000;
		12'd0747: rd_data_0 <= 24'hff0000;
		12'd0748: rd_data_0 <= 24'hff0000;
		12'd0749: rd_data_0 <= 24'hff0000;
		12'd0750: rd_data_0 <= 24'hff0000;
		12'd0751: rd_data_0 <= 24'hff0000;
		12'd0752: rd_data_0 <= 24'h0000ff;
		12'd0753: rd_data_0 <= 24'h0000ff;
		12'd0754: rd_data_0 <= 24'h0000ff;
		12'd0755: rd_data_0 <= 24'h0000ff;
		12'd0756: rd_data_0 <= 24'h0000ff;
		12'd0757: rd_data_0 <= 24'h0000ff;
		12'd0758: rd_data_0 <= 24'h0000ff;
		12'd0759: rd_data_0 <= 24'h0000ff;
		12'd0760: rd_data_0 <= 24'h000000;
		12'd0761: rd_data_0 <= 24'h000000;
		12'd0762: rd_data_0 <= 24'h000000;
		12'd0763: rd_data_0 <= 24'h000000;
		12'd0764: rd_data_0 <= 24'h000000;
		12'd0765: rd_data_0 <= 24'h000000;
		12'd0766: rd_data_0 <= 24'h000000;
		12'd0767: rd_data_0 <= 24'h000000;
		12'd0768: rd_data_0 <= 24'hffffff;
		12'd0769: rd_data_0 <= 24'hffffff;
		12'd0770: rd_data_0 <= 24'hffffff;
		12'd0771: rd_data_0 <= 24'hffffff;
		12'd0772: rd_data_0 <= 24'hffffff;
		12'd0773: rd_data_0 <= 24'hffffff;
		12'd0774: rd_data_0 <= 24'hffffff;
		12'd0775: rd_data_0 <= 24'hffffff;
		12'd0776: rd_data_0 <= 24'hffff00;
		12'd0777: rd_data_0 <= 24'hffff00;
		12'd0778: rd_data_0 <= 24'hffff00;
		12'd0779: rd_data_0 <= 24'hffff00;
		12'd0780: rd_data_0 <= 24'hffff00;
		12'd0781: rd_data_0 <= 24'hffff00;
		12'd0782: rd_data_0 <= 24'hffff00;
		12'd0783: rd_data_0 <= 24'hffff00;
		12'd0784: rd_data_0 <= 24'h00ffff;
		12'd0785: rd_data_0 <= 24'h00ffff;
		12'd0786: rd_data_0 <= 24'h00ffff;
		12'd0787: rd_data_0 <= 24'h00ffff;
		12'd0788: rd_data_0 <= 24'h00ffff;
		12'd0789: rd_data_0 <= 24'h00ffff;
		12'd0790: rd_data_0 <= 24'h00ffff;
		12'd0791: rd_data_0 <= 24'h00ffff;
		12'd0792: rd_data_0 <= 24'h00ff00;
		12'd0793: rd_data_0 <= 24'h00ff00;
		12'd0794: rd_data_0 <= 24'h00ff00;
		12'd0795: rd_data_0 <= 24'h00ff00;
		12'd0796: rd_data_0 <= 24'h00ff00;
		12'd0797: rd_data_0 <= 24'h00ff00;
		12'd0798: rd_data_0 <= 24'h00ff00;
		12'd0799: rd_data_0 <= 24'h00ff00;
		12'd0800: rd_data_0 <= 24'hff00ff;
		12'd0801: rd_data_0 <= 24'hff00ff;
		12'd0802: rd_data_0 <= 24'hff00ff;
		12'd0803: rd_data_0 <= 24'hff00ff;
		12'd0804: rd_data_0 <= 24'hff00ff;
		12'd0805: rd_data_0 <= 24'hff00ff;
		12'd0806: rd_data_0 <= 24'hff00ff;
		12'd0807: rd_data_0 <= 24'hff00ff;
		12'd0808: rd_data_0 <= 24'hff0000;
		12'd0809: rd_data_0 <= 24'hff0000;
		12'd0810: rd_data_0 <= 24'hff0000;
		12'd0811: rd_data_0 <= 24'hff0000;
		12'd0812: rd_data_0 <= 24'hff0000;
		12'd0813: rd_data_0 <= 24'hff0000;
		12'd0814: rd_data_0 <= 24'hff0000;
		12'd0815: rd_data_0 <= 24'hff0000;
		12'd0816: rd_data_0 <= 24'h0000ff;
		12'd0817: rd_data_0 <= 24'h0000ff;
		12'd0818: rd_data_0 <= 24'h0000ff;
		12'd0819: rd_data_0 <= 24'h0000ff;
		12'd0820: rd_data_0 <= 24'h0000ff;
		12'd0821: rd_data_0 <= 24'h0000ff;
		12'd0822: rd_data_0 <= 24'h0000ff;
		12'd0823: rd_data_0 <= 24'h0000ff;
		12'd0824: rd_data_0 <= 24'h000000;
		12'd0825: rd_data_0 <= 24'h000000;
		12'd0826: rd_data_0 <= 24'h000000;
		12'd0827: rd_data_0 <= 24'h000000;
		12'd0828: rd_data_0 <= 24'h000000;
		12'd0829: rd_data_0 <= 24'h000000;
		12'd0830: rd_data_0 <= 24'h000000;
		12'd0831: rd_data_0 <= 24'h000000;
		12'd0832: rd_data_0 <= 24'hffffff;
		12'd0833: rd_data_0 <= 24'hffffff;
		12'd0834: rd_data_0 <= 24'hffffff;
		12'd0835: rd_data_0 <= 24'hffffff;
		12'd0836: rd_data_0 <= 24'hffffff;
		12'd0837: rd_data_0 <= 24'hffffff;
		12'd0838: rd_data_0 <= 24'hffffff;
		12'd0839: rd_data_0 <= 24'hffffff;
		12'd0840: rd_data_0 <= 24'hffff00;
		12'd0841: rd_data_0 <= 24'hffff00;
		12'd0842: rd_data_0 <= 24'hffff00;
		12'd0843: rd_data_0 <= 24'hffff00;
		12'd0844: rd_data_0 <= 24'hffff00;
		12'd0845: rd_data_0 <= 24'hffff00;
		12'd0846: rd_data_0 <= 24'hffff00;
		12'd0847: rd_data_0 <= 24'hffff00;
		12'd0848: rd_data_0 <= 24'h00ffff;
		12'd0849: rd_data_0 <= 24'h00ffff;
		12'd0850: rd_data_0 <= 24'h00ffff;
		12'd0851: rd_data_0 <= 24'h00ffff;
		12'd0852: rd_data_0 <= 24'h00ffff;
		12'd0853: rd_data_0 <= 24'h00ffff;
		12'd0854: rd_data_0 <= 24'h00ffff;
		12'd0855: rd_data_0 <= 24'h00ffff;
		12'd0856: rd_data_0 <= 24'h00ff00;
		12'd0857: rd_data_0 <= 24'h00ff00;
		12'd0858: rd_data_0 <= 24'h00ff00;
		12'd0859: rd_data_0 <= 24'h00ff00;
		12'd0860: rd_data_0 <= 24'h00ff00;
		12'd0861: rd_data_0 <= 24'h00ff00;
		12'd0862: rd_data_0 <= 24'h00ff00;
		12'd0863: rd_data_0 <= 24'h00ff00;
		12'd0864: rd_data_0 <= 24'hff00ff;
		12'd0865: rd_data_0 <= 24'hff00ff;
		12'd0866: rd_data_0 <= 24'hff00ff;
		12'd0867: rd_data_0 <= 24'hff00ff;
		12'd0868: rd_data_0 <= 24'hff00ff;
		12'd0869: rd_data_0 <= 24'hff00ff;
		12'd0870: rd_data_0 <= 24'hff00ff;
		12'd0871: rd_data_0 <= 24'hff00ff;
		12'd0872: rd_data_0 <= 24'hff0000;
		12'd0873: rd_data_0 <= 24'hff0000;
		12'd0874: rd_data_0 <= 24'hff0000;
		12'd0875: rd_data_0 <= 24'hff0000;
		12'd0876: rd_data_0 <= 24'hff0000;
		12'd0877: rd_data_0 <= 24'hff0000;
		12'd0878: rd_data_0 <= 24'hff0000;
		12'd0879: rd_data_0 <= 24'hff0000;
		12'd0880: rd_data_0 <= 24'h0000ff;
		12'd0881: rd_data_0 <= 24'h0000ff;
		12'd0882: rd_data_0 <= 24'h0000ff;
		12'd0883: rd_data_0 <= 24'h0000ff;
		12'd0884: rd_data_0 <= 24'h0000ff;
		12'd0885: rd_data_0 <= 24'h0000ff;
		12'd0886: rd_data_0 <= 24'h0000ff;
		12'd0887: rd_data_0 <= 24'h0000ff;
		12'd0888: rd_data_0 <= 24'h000000;
		12'd0889: rd_data_0 <= 24'h000000;
		12'd0890: rd_data_0 <= 24'h000000;
		12'd0891: rd_data_0 <= 24'h000000;
		12'd0892: rd_data_0 <= 24'h000000;
		12'd0893: rd_data_0 <= 24'h000000;
		12'd0894: rd_data_0 <= 24'h000000;
		12'd0895: rd_data_0 <= 24'h000000;
		12'd0896: rd_data_0 <= 24'hffffff;
		12'd0897: rd_data_0 <= 24'hffffff;
		12'd0898: rd_data_0 <= 24'hffffff;
		12'd0899: rd_data_0 <= 24'hffffff;
		12'd0900: rd_data_0 <= 24'hffffff;
		12'd0901: rd_data_0 <= 24'hffffff;
		12'd0902: rd_data_0 <= 24'hffffff;
		12'd0903: rd_data_0 <= 24'hffffff;
		12'd0904: rd_data_0 <= 24'hffff00;
		12'd0905: rd_data_0 <= 24'hffff00;
		12'd0906: rd_data_0 <= 24'hffff00;
		12'd0907: rd_data_0 <= 24'hffff00;
		12'd0908: rd_data_0 <= 24'hffff00;
		12'd0909: rd_data_0 <= 24'hffff00;
		12'd0910: rd_data_0 <= 24'hffff00;
		12'd0911: rd_data_0 <= 24'hffff00;
		12'd0912: rd_data_0 <= 24'h00ffff;
		12'd0913: rd_data_0 <= 24'h00ffff;
		12'd0914: rd_data_0 <= 24'h00ffff;
		12'd0915: rd_data_0 <= 24'h00ffff;
		12'd0916: rd_data_0 <= 24'h00ffff;
		12'd0917: rd_data_0 <= 24'h00ffff;
		12'd0918: rd_data_0 <= 24'h00ffff;
		12'd0919: rd_data_0 <= 24'h00ffff;
		12'd0920: rd_data_0 <= 24'h00ff00;
		12'd0921: rd_data_0 <= 24'h00ff00;
		12'd0922: rd_data_0 <= 24'h00ff00;
		12'd0923: rd_data_0 <= 24'h00ff00;
		12'd0924: rd_data_0 <= 24'h00ff00;
		12'd0925: rd_data_0 <= 24'h00ff00;
		12'd0926: rd_data_0 <= 24'h00ff00;
		12'd0927: rd_data_0 <= 24'h00ff00;
		12'd0928: rd_data_0 <= 24'hff00ff;
		12'd0929: rd_data_0 <= 24'hff00ff;
		12'd0930: rd_data_0 <= 24'hff00ff;
		12'd0931: rd_data_0 <= 24'hff00ff;
		12'd0932: rd_data_0 <= 24'hff00ff;
		12'd0933: rd_data_0 <= 24'hff00ff;
		12'd0934: rd_data_0 <= 24'hff00ff;
		12'd0935: rd_data_0 <= 24'hff00ff;
		12'd0936: rd_data_0 <= 24'hff0000;
		12'd0937: rd_data_0 <= 24'hff0000;
		12'd0938: rd_data_0 <= 24'hff0000;
		12'd0939: rd_data_0 <= 24'hff0000;
		12'd0940: rd_data_0 <= 24'hff0000;
		12'd0941: rd_data_0 <= 24'hff0000;
		12'd0942: rd_data_0 <= 24'hff0000;
		12'd0943: rd_data_0 <= 24'hff0000;
		12'd0944: rd_data_0 <= 24'h0000ff;
		12'd0945: rd_data_0 <= 24'h0000ff;
		12'd0946: rd_data_0 <= 24'h0000ff;
		12'd0947: rd_data_0 <= 24'h0000ff;
		12'd0948: rd_data_0 <= 24'h0000ff;
		12'd0949: rd_data_0 <= 24'h0000ff;
		12'd0950: rd_data_0 <= 24'h0000ff;
		12'd0951: rd_data_0 <= 24'h0000ff;
		12'd0952: rd_data_0 <= 24'h000000;
		12'd0953: rd_data_0 <= 24'h000000;
		12'd0954: rd_data_0 <= 24'h000000;
		12'd0955: rd_data_0 <= 24'h000000;
		12'd0956: rd_data_0 <= 24'h000000;
		12'd0957: rd_data_0 <= 24'h000000;
		12'd0958: rd_data_0 <= 24'h000000;
		12'd0959: rd_data_0 <= 24'h000000;
		12'd0960: rd_data_0 <= 24'hffffff;
		12'd0961: rd_data_0 <= 24'hffffff;
		12'd0962: rd_data_0 <= 24'hffffff;
		12'd0963: rd_data_0 <= 24'hffffff;
		12'd0964: rd_data_0 <= 24'hffffff;
		12'd0965: rd_data_0 <= 24'hffffff;
		12'd0966: rd_data_0 <= 24'hffffff;
		12'd0967: rd_data_0 <= 24'hffffff;
		12'd0968: rd_data_0 <= 24'hffff00;
		12'd0969: rd_data_0 <= 24'hffff00;
		12'd0970: rd_data_0 <= 24'hffff00;
		12'd0971: rd_data_0 <= 24'hffff00;
		12'd0972: rd_data_0 <= 24'hffff00;
		12'd0973: rd_data_0 <= 24'hffff00;
		12'd0974: rd_data_0 <= 24'hffff00;
		12'd0975: rd_data_0 <= 24'hffff00;
		12'd0976: rd_data_0 <= 24'h00ffff;
		12'd0977: rd_data_0 <= 24'h00ffff;
		12'd0978: rd_data_0 <= 24'h00ffff;
		12'd0979: rd_data_0 <= 24'h00ffff;
		12'd0980: rd_data_0 <= 24'h00ffff;
		12'd0981: rd_data_0 <= 24'h00ffff;
		12'd0982: rd_data_0 <= 24'h00ffff;
		12'd0983: rd_data_0 <= 24'h00ffff;
		12'd0984: rd_data_0 <= 24'h00ff00;
		12'd0985: rd_data_0 <= 24'h00ff00;
		12'd0986: rd_data_0 <= 24'h00ff00;
		12'd0987: rd_data_0 <= 24'h00ff00;
		12'd0988: rd_data_0 <= 24'h00ff00;
		12'd0989: rd_data_0 <= 24'h00ff00;
		12'd0990: rd_data_0 <= 24'h00ff00;
		12'd0991: rd_data_0 <= 24'h00ff00;
		12'd0992: rd_data_0 <= 24'hff00ff;
		12'd0993: rd_data_0 <= 24'hff00ff;
		12'd0994: rd_data_0 <= 24'hff00ff;
		12'd0995: rd_data_0 <= 24'hff00ff;
		12'd0996: rd_data_0 <= 24'hff00ff;
		12'd0997: rd_data_0 <= 24'hff00ff;
		12'd0998: rd_data_0 <= 24'hff00ff;
		12'd0999: rd_data_0 <= 24'hff00ff;
		12'd1000: rd_data_0 <= 24'hff0000;
		12'd1001: rd_data_0 <= 24'hff0000;
		12'd1002: rd_data_0 <= 24'hff0000;
		12'd1003: rd_data_0 <= 24'hff0000;
		12'd1004: rd_data_0 <= 24'hff0000;
		12'd1005: rd_data_0 <= 24'hff0000;
		12'd1006: rd_data_0 <= 24'hff0000;
		12'd1007: rd_data_0 <= 24'hff0000;
		12'd1008: rd_data_0 <= 24'h0000ff;
		12'd1009: rd_data_0 <= 24'h0000ff;
		12'd1010: rd_data_0 <= 24'h0000ff;
		12'd1011: rd_data_0 <= 24'h0000ff;
		12'd1012: rd_data_0 <= 24'h0000ff;
		12'd1013: rd_data_0 <= 24'h0000ff;
		12'd1014: rd_data_0 <= 24'h0000ff;
		12'd1015: rd_data_0 <= 24'h0000ff;
		12'd1016: rd_data_0 <= 24'h000000;
		12'd1017: rd_data_0 <= 24'h000000;
		12'd1018: rd_data_0 <= 24'h000000;
		12'd1019: rd_data_0 <= 24'h000000;
		12'd1020: rd_data_0 <= 24'h000000;
		12'd1021: rd_data_0 <= 24'h000000;
		12'd1022: rd_data_0 <= 24'h000000;
		12'd1023: rd_data_0 <= 24'h000000;
		12'd1024: rd_data_0 <= 24'hffffff;
		12'd1025: rd_data_0 <= 24'hffffff;
		12'd1026: rd_data_0 <= 24'hffffff;
		12'd1027: rd_data_0 <= 24'hffffff;
		12'd1028: rd_data_0 <= 24'hffffff;
		12'd1029: rd_data_0 <= 24'hffffff;
		12'd1030: rd_data_0 <= 24'hffffff;
		12'd1031: rd_data_0 <= 24'hffffff;
		12'd1032: rd_data_0 <= 24'hffff00;
		12'd1033: rd_data_0 <= 24'hffff00;
		12'd1034: rd_data_0 <= 24'hffff00;
		12'd1035: rd_data_0 <= 24'hffff00;
		12'd1036: rd_data_0 <= 24'hffff00;
		12'd1037: rd_data_0 <= 24'hffff00;
		12'd1038: rd_data_0 <= 24'hffff00;
		12'd1039: rd_data_0 <= 24'hffff00;
		12'd1040: rd_data_0 <= 24'h00ffff;
		12'd1041: rd_data_0 <= 24'h00ffff;
		12'd1042: rd_data_0 <= 24'h00ffff;
		12'd1043: rd_data_0 <= 24'h00ffff;
		12'd1044: rd_data_0 <= 24'h00ffff;
		12'd1045: rd_data_0 <= 24'h00ffff;
		12'd1046: rd_data_0 <= 24'h00ffff;
		12'd1047: rd_data_0 <= 24'h00ffff;
		12'd1048: rd_data_0 <= 24'h00ff00;
		12'd1049: rd_data_0 <= 24'h00ff00;
		12'd1050: rd_data_0 <= 24'h00ff00;
		12'd1051: rd_data_0 <= 24'h00ff00;
		12'd1052: rd_data_0 <= 24'h00ff00;
		12'd1053: rd_data_0 <= 24'h00ff00;
		12'd1054: rd_data_0 <= 24'h00ff00;
		12'd1055: rd_data_0 <= 24'h00ff00;
		12'd1056: rd_data_0 <= 24'hff00ff;
		12'd1057: rd_data_0 <= 24'hff00ff;
		12'd1058: rd_data_0 <= 24'hff00ff;
		12'd1059: rd_data_0 <= 24'hff00ff;
		12'd1060: rd_data_0 <= 24'hff00ff;
		12'd1061: rd_data_0 <= 24'hff00ff;
		12'd1062: rd_data_0 <= 24'hff00ff;
		12'd1063: rd_data_0 <= 24'hff00ff;
		12'd1064: rd_data_0 <= 24'hff0000;
		12'd1065: rd_data_0 <= 24'hff0000;
		12'd1066: rd_data_0 <= 24'hff0000;
		12'd1067: rd_data_0 <= 24'hff0000;
		12'd1068: rd_data_0 <= 24'hff0000;
		12'd1069: rd_data_0 <= 24'hff0000;
		12'd1070: rd_data_0 <= 24'hff0000;
		12'd1071: rd_data_0 <= 24'hff0000;
		12'd1072: rd_data_0 <= 24'h0000ff;
		12'd1073: rd_data_0 <= 24'h0000ff;
		12'd1074: rd_data_0 <= 24'h0000ff;
		12'd1075: rd_data_0 <= 24'h0000ff;
		12'd1076: rd_data_0 <= 24'h0000ff;
		12'd1077: rd_data_0 <= 24'h0000ff;
		12'd1078: rd_data_0 <= 24'h0000ff;
		12'd1079: rd_data_0 <= 24'h0000ff;
		12'd1080: rd_data_0 <= 24'h000000;
		12'd1081: rd_data_0 <= 24'h000000;
		12'd1082: rd_data_0 <= 24'h000000;
		12'd1083: rd_data_0 <= 24'h000000;
		12'd1084: rd_data_0 <= 24'h000000;
		12'd1085: rd_data_0 <= 24'h000000;
		12'd1086: rd_data_0 <= 24'h000000;
		12'd1087: rd_data_0 <= 24'h000000;
		12'd1088: rd_data_0 <= 24'hffffff;
		12'd1089: rd_data_0 <= 24'hffffff;
		12'd1090: rd_data_0 <= 24'hffffff;
		12'd1091: rd_data_0 <= 24'hffffff;
		12'd1092: rd_data_0 <= 24'hffffff;
		12'd1093: rd_data_0 <= 24'hffffff;
		12'd1094: rd_data_0 <= 24'hffffff;
		12'd1095: rd_data_0 <= 24'hffffff;
		12'd1096: rd_data_0 <= 24'hffff00;
		12'd1097: rd_data_0 <= 24'hffff00;
		12'd1098: rd_data_0 <= 24'hffff00;
		12'd1099: rd_data_0 <= 24'hffff00;
		12'd1100: rd_data_0 <= 24'hffff00;
		12'd1101: rd_data_0 <= 24'hffff00;
		12'd1102: rd_data_0 <= 24'hffff00;
		12'd1103: rd_data_0 <= 24'hffff00;
		12'd1104: rd_data_0 <= 24'h00ffff;
		12'd1105: rd_data_0 <= 24'h00ffff;
		12'd1106: rd_data_0 <= 24'h00ffff;
		12'd1107: rd_data_0 <= 24'h00ffff;
		12'd1108: rd_data_0 <= 24'h00ffff;
		12'd1109: rd_data_0 <= 24'h00ffff;
		12'd1110: rd_data_0 <= 24'h00ffff;
		12'd1111: rd_data_0 <= 24'h00ffff;
		12'd1112: rd_data_0 <= 24'h00ff00;
		12'd1113: rd_data_0 <= 24'h00ff00;
		12'd1114: rd_data_0 <= 24'h00ff00;
		12'd1115: rd_data_0 <= 24'h00ff00;
		12'd1116: rd_data_0 <= 24'h00ff00;
		12'd1117: rd_data_0 <= 24'h00ff00;
		12'd1118: rd_data_0 <= 24'h00ff00;
		12'd1119: rd_data_0 <= 24'h00ff00;
		12'd1120: rd_data_0 <= 24'hff00ff;
		12'd1121: rd_data_0 <= 24'hff00ff;
		12'd1122: rd_data_0 <= 24'hff00ff;
		12'd1123: rd_data_0 <= 24'hff00ff;
		12'd1124: rd_data_0 <= 24'hff00ff;
		12'd1125: rd_data_0 <= 24'hff00ff;
		12'd1126: rd_data_0 <= 24'hff00ff;
		12'd1127: rd_data_0 <= 24'hff00ff;
		12'd1128: rd_data_0 <= 24'hff0000;
		12'd1129: rd_data_0 <= 24'hff0000;
		12'd1130: rd_data_0 <= 24'hff0000;
		12'd1131: rd_data_0 <= 24'hff0000;
		12'd1132: rd_data_0 <= 24'hff0000;
		12'd1133: rd_data_0 <= 24'hff0000;
		12'd1134: rd_data_0 <= 24'hff0000;
		12'd1135: rd_data_0 <= 24'hff0000;
		12'd1136: rd_data_0 <= 24'h0000ff;
		12'd1137: rd_data_0 <= 24'h0000ff;
		12'd1138: rd_data_0 <= 24'h0000ff;
		12'd1139: rd_data_0 <= 24'h0000ff;
		12'd1140: rd_data_0 <= 24'h0000ff;
		12'd1141: rd_data_0 <= 24'h0000ff;
		12'd1142: rd_data_0 <= 24'h0000ff;
		12'd1143: rd_data_0 <= 24'h0000ff;
		12'd1144: rd_data_0 <= 24'h000000;
		12'd1145: rd_data_0 <= 24'h000000;
		12'd1146: rd_data_0 <= 24'h000000;
		12'd1147: rd_data_0 <= 24'h000000;
		12'd1148: rd_data_0 <= 24'h000000;
		12'd1149: rd_data_0 <= 24'h000000;
		12'd1150: rd_data_0 <= 24'h000000;
		12'd1151: rd_data_0 <= 24'h000000;
		12'd1152: rd_data_0 <= 24'hffffff;
		12'd1153: rd_data_0 <= 24'hffffff;
		12'd1154: rd_data_0 <= 24'hffffff;
		12'd1155: rd_data_0 <= 24'hffffff;
		12'd1156: rd_data_0 <= 24'hffffff;
		12'd1157: rd_data_0 <= 24'hffffff;
		12'd1158: rd_data_0 <= 24'hffffff;
		12'd1159: rd_data_0 <= 24'hffffff;
		12'd1160: rd_data_0 <= 24'hffff00;
		12'd1161: rd_data_0 <= 24'hffff00;
		12'd1162: rd_data_0 <= 24'hffff00;
		12'd1163: rd_data_0 <= 24'hffff00;
		12'd1164: rd_data_0 <= 24'hffff00;
		12'd1165: rd_data_0 <= 24'hffff00;
		12'd1166: rd_data_0 <= 24'hffff00;
		12'd1167: rd_data_0 <= 24'hffff00;
		12'd1168: rd_data_0 <= 24'h00ffff;
		12'd1169: rd_data_0 <= 24'h00ffff;
		12'd1170: rd_data_0 <= 24'h00ffff;
		12'd1171: rd_data_0 <= 24'h00ffff;
		12'd1172: rd_data_0 <= 24'h00ffff;
		12'd1173: rd_data_0 <= 24'h00ffff;
		12'd1174: rd_data_0 <= 24'h00ffff;
		12'd1175: rd_data_0 <= 24'h00ffff;
		12'd1176: rd_data_0 <= 24'h00ff00;
		12'd1177: rd_data_0 <= 24'h00ff00;
		12'd1178: rd_data_0 <= 24'h00ff00;
		12'd1179: rd_data_0 <= 24'h00ff00;
		12'd1180: rd_data_0 <= 24'h00ff00;
		12'd1181: rd_data_0 <= 24'h00ff00;
		12'd1182: rd_data_0 <= 24'h00ff00;
		12'd1183: rd_data_0 <= 24'h00ff00;
		12'd1184: rd_data_0 <= 24'hff00ff;
		12'd1185: rd_data_0 <= 24'hff00ff;
		12'd1186: rd_data_0 <= 24'hff00ff;
		12'd1187: rd_data_0 <= 24'hff00ff;
		12'd1188: rd_data_0 <= 24'hff00ff;
		12'd1189: rd_data_0 <= 24'hff00ff;
		12'd1190: rd_data_0 <= 24'hff00ff;
		12'd1191: rd_data_0 <= 24'hff00ff;
		12'd1192: rd_data_0 <= 24'hff0000;
		12'd1193: rd_data_0 <= 24'hff0000;
		12'd1194: rd_data_0 <= 24'hff0000;
		12'd1195: rd_data_0 <= 24'hff0000;
		12'd1196: rd_data_0 <= 24'hff0000;
		12'd1197: rd_data_0 <= 24'hff0000;
		12'd1198: rd_data_0 <= 24'hff0000;
		12'd1199: rd_data_0 <= 24'hff0000;
		12'd1200: rd_data_0 <= 24'h0000ff;
		12'd1201: rd_data_0 <= 24'h0000ff;
		12'd1202: rd_data_0 <= 24'h0000ff;
		12'd1203: rd_data_0 <= 24'h0000ff;
		12'd1204: rd_data_0 <= 24'h0000ff;
		12'd1205: rd_data_0 <= 24'h0000ff;
		12'd1206: rd_data_0 <= 24'h0000ff;
		12'd1207: rd_data_0 <= 24'h0000ff;
		12'd1208: rd_data_0 <= 24'h000000;
		12'd1209: rd_data_0 <= 24'h000000;
		12'd1210: rd_data_0 <= 24'h000000;
		12'd1211: rd_data_0 <= 24'h000000;
		12'd1212: rd_data_0 <= 24'h000000;
		12'd1213: rd_data_0 <= 24'h000000;
		12'd1214: rd_data_0 <= 24'h000000;
		12'd1215: rd_data_0 <= 24'h000000;
		12'd1216: rd_data_0 <= 24'hffffff;
		12'd1217: rd_data_0 <= 24'hffffff;
		12'd1218: rd_data_0 <= 24'hffffff;
		12'd1219: rd_data_0 <= 24'hffffff;
		12'd1220: rd_data_0 <= 24'hffffff;
		12'd1221: rd_data_0 <= 24'hffffff;
		12'd1222: rd_data_0 <= 24'hffffff;
		12'd1223: rd_data_0 <= 24'hffffff;
		12'd1224: rd_data_0 <= 24'hffff00;
		12'd1225: rd_data_0 <= 24'hffff00;
		12'd1226: rd_data_0 <= 24'hffff00;
		12'd1227: rd_data_0 <= 24'hffff00;
		12'd1228: rd_data_0 <= 24'hffff00;
		12'd1229: rd_data_0 <= 24'hffff00;
		12'd1230: rd_data_0 <= 24'hffff00;
		12'd1231: rd_data_0 <= 24'hffff00;
		12'd1232: rd_data_0 <= 24'h00ffff;
		12'd1233: rd_data_0 <= 24'h00ffff;
		12'd1234: rd_data_0 <= 24'h00ffff;
		12'd1235: rd_data_0 <= 24'h00ffff;
		12'd1236: rd_data_0 <= 24'h00ffff;
		12'd1237: rd_data_0 <= 24'h00ffff;
		12'd1238: rd_data_0 <= 24'h00ffff;
		12'd1239: rd_data_0 <= 24'h00ffff;
		12'd1240: rd_data_0 <= 24'h00ff00;
		12'd1241: rd_data_0 <= 24'h00ff00;
		12'd1242: rd_data_0 <= 24'h00ff00;
		12'd1243: rd_data_0 <= 24'h00ff00;
		12'd1244: rd_data_0 <= 24'h00ff00;
		12'd1245: rd_data_0 <= 24'h00ff00;
		12'd1246: rd_data_0 <= 24'h00ff00;
		12'd1247: rd_data_0 <= 24'h00ff00;
		12'd1248: rd_data_0 <= 24'hff00ff;
		12'd1249: rd_data_0 <= 24'hff00ff;
		12'd1250: rd_data_0 <= 24'hff00ff;
		12'd1251: rd_data_0 <= 24'hff00ff;
		12'd1252: rd_data_0 <= 24'hff00ff;
		12'd1253: rd_data_0 <= 24'hff00ff;
		12'd1254: rd_data_0 <= 24'hff00ff;
		12'd1255: rd_data_0 <= 24'hff00ff;
		12'd1256: rd_data_0 <= 24'hff0000;
		12'd1257: rd_data_0 <= 24'hff0000;
		12'd1258: rd_data_0 <= 24'hff0000;
		12'd1259: rd_data_0 <= 24'hff0000;
		12'd1260: rd_data_0 <= 24'hff0000;
		12'd1261: rd_data_0 <= 24'hff0000;
		12'd1262: rd_data_0 <= 24'hff0000;
		12'd1263: rd_data_0 <= 24'hff0000;
		12'd1264: rd_data_0 <= 24'h0000ff;
		12'd1265: rd_data_0 <= 24'h0000ff;
		12'd1266: rd_data_0 <= 24'h0000ff;
		12'd1267: rd_data_0 <= 24'h0000ff;
		12'd1268: rd_data_0 <= 24'h0000ff;
		12'd1269: rd_data_0 <= 24'h0000ff;
		12'd1270: rd_data_0 <= 24'h0000ff;
		12'd1271: rd_data_0 <= 24'h0000ff;
		12'd1272: rd_data_0 <= 24'h000000;
		12'd1273: rd_data_0 <= 24'h000000;
		12'd1274: rd_data_0 <= 24'h000000;
		12'd1275: rd_data_0 <= 24'h000000;
		12'd1276: rd_data_0 <= 24'h000000;
		12'd1277: rd_data_0 <= 24'h000000;
		12'd1278: rd_data_0 <= 24'h000000;
		12'd1279: rd_data_0 <= 24'h000000;
		12'd1280: rd_data_0 <= 24'hffffff;
		12'd1281: rd_data_0 <= 24'hffffff;
		12'd1282: rd_data_0 <= 24'hffffff;
		12'd1283: rd_data_0 <= 24'hffffff;
		12'd1284: rd_data_0 <= 24'hffffff;
		12'd1285: rd_data_0 <= 24'hffffff;
		12'd1286: rd_data_0 <= 24'hffffff;
		12'd1287: rd_data_0 <= 24'hffffff;
		12'd1288: rd_data_0 <= 24'hffff00;
		12'd1289: rd_data_0 <= 24'hffff00;
		12'd1290: rd_data_0 <= 24'hffff00;
		12'd1291: rd_data_0 <= 24'hffff00;
		12'd1292: rd_data_0 <= 24'hffff00;
		12'd1293: rd_data_0 <= 24'hffff00;
		12'd1294: rd_data_0 <= 24'hffff00;
		12'd1295: rd_data_0 <= 24'hffff00;
		12'd1296: rd_data_0 <= 24'h00ffff;
		12'd1297: rd_data_0 <= 24'h00ffff;
		12'd1298: rd_data_0 <= 24'h00ffff;
		12'd1299: rd_data_0 <= 24'h00ffff;
		12'd1300: rd_data_0 <= 24'h00ffff;
		12'd1301: rd_data_0 <= 24'h00ffff;
		12'd1302: rd_data_0 <= 24'h00ffff;
		12'd1303: rd_data_0 <= 24'h00ffff;
		12'd1304: rd_data_0 <= 24'h00ff00;
		12'd1305: rd_data_0 <= 24'h00ff00;
		12'd1306: rd_data_0 <= 24'h00ff00;
		12'd1307: rd_data_0 <= 24'h00ff00;
		12'd1308: rd_data_0 <= 24'h00ff00;
		12'd1309: rd_data_0 <= 24'h00ff00;
		12'd1310: rd_data_0 <= 24'h00ff00;
		12'd1311: rd_data_0 <= 24'h00ff00;
		12'd1312: rd_data_0 <= 24'hff00ff;
		12'd1313: rd_data_0 <= 24'hff00ff;
		12'd1314: rd_data_0 <= 24'hff00ff;
		12'd1315: rd_data_0 <= 24'hff00ff;
		12'd1316: rd_data_0 <= 24'hff00ff;
		12'd1317: rd_data_0 <= 24'hff00ff;
		12'd1318: rd_data_0 <= 24'hff00ff;
		12'd1319: rd_data_0 <= 24'hff00ff;
		12'd1320: rd_data_0 <= 24'hff0000;
		12'd1321: rd_data_0 <= 24'hff0000;
		12'd1322: rd_data_0 <= 24'hff0000;
		12'd1323: rd_data_0 <= 24'hff0000;
		12'd1324: rd_data_0 <= 24'hff0000;
		12'd1325: rd_data_0 <= 24'hff0000;
		12'd1326: rd_data_0 <= 24'hff0000;
		12'd1327: rd_data_0 <= 24'hff0000;
		12'd1328: rd_data_0 <= 24'h0000ff;
		12'd1329: rd_data_0 <= 24'h0000ff;
		12'd1330: rd_data_0 <= 24'h0000ff;
		12'd1331: rd_data_0 <= 24'h0000ff;
		12'd1332: rd_data_0 <= 24'h0000ff;
		12'd1333: rd_data_0 <= 24'h0000ff;
		12'd1334: rd_data_0 <= 24'h0000ff;
		12'd1335: rd_data_0 <= 24'h0000ff;
		12'd1336: rd_data_0 <= 24'h000000;
		12'd1337: rd_data_0 <= 24'h000000;
		12'd1338: rd_data_0 <= 24'h000000;
		12'd1339: rd_data_0 <= 24'h000000;
		12'd1340: rd_data_0 <= 24'h000000;
		12'd1341: rd_data_0 <= 24'h000000;
		12'd1342: rd_data_0 <= 24'h000000;
		12'd1343: rd_data_0 <= 24'h000000;
		12'd1344: rd_data_0 <= 24'hffffff;
		12'd1345: rd_data_0 <= 24'hffffff;
		12'd1346: rd_data_0 <= 24'hffffff;
		12'd1347: rd_data_0 <= 24'hffffff;
		12'd1348: rd_data_0 <= 24'hffffff;
		12'd1349: rd_data_0 <= 24'hffffff;
		12'd1350: rd_data_0 <= 24'hffffff;
		12'd1351: rd_data_0 <= 24'hffffff;
		12'd1352: rd_data_0 <= 24'hffff00;
		12'd1353: rd_data_0 <= 24'hffff00;
		12'd1354: rd_data_0 <= 24'hffff00;
		12'd1355: rd_data_0 <= 24'hffff00;
		12'd1356: rd_data_0 <= 24'hffff00;
		12'd1357: rd_data_0 <= 24'hffff00;
		12'd1358: rd_data_0 <= 24'hffff00;
		12'd1359: rd_data_0 <= 24'hffff00;
		12'd1360: rd_data_0 <= 24'h00ffff;
		12'd1361: rd_data_0 <= 24'h00ffff;
		12'd1362: rd_data_0 <= 24'h00ffff;
		12'd1363: rd_data_0 <= 24'h00ffff;
		12'd1364: rd_data_0 <= 24'h00ffff;
		12'd1365: rd_data_0 <= 24'h00ffff;
		12'd1366: rd_data_0 <= 24'h00ffff;
		12'd1367: rd_data_0 <= 24'h00ffff;
		12'd1368: rd_data_0 <= 24'h00ff00;
		12'd1369: rd_data_0 <= 24'h00ff00;
		12'd1370: rd_data_0 <= 24'h00ff00;
		12'd1371: rd_data_0 <= 24'h00ff00;
		12'd1372: rd_data_0 <= 24'h00ff00;
		12'd1373: rd_data_0 <= 24'h00ff00;
		12'd1374: rd_data_0 <= 24'h00ff00;
		12'd1375: rd_data_0 <= 24'h00ff00;
		12'd1376: rd_data_0 <= 24'hff00ff;
		12'd1377: rd_data_0 <= 24'hff00ff;
		12'd1378: rd_data_0 <= 24'hff00ff;
		12'd1379: rd_data_0 <= 24'hff00ff;
		12'd1380: rd_data_0 <= 24'hff00ff;
		12'd1381: rd_data_0 <= 24'hff00ff;
		12'd1382: rd_data_0 <= 24'hff00ff;
		12'd1383: rd_data_0 <= 24'hff00ff;
		12'd1384: rd_data_0 <= 24'hff0000;
		12'd1385: rd_data_0 <= 24'hff0000;
		12'd1386: rd_data_0 <= 24'hff0000;
		12'd1387: rd_data_0 <= 24'hff0000;
		12'd1388: rd_data_0 <= 24'hff0000;
		12'd1389: rd_data_0 <= 24'hff0000;
		12'd1390: rd_data_0 <= 24'hff0000;
		12'd1391: rd_data_0 <= 24'hff0000;
		12'd1392: rd_data_0 <= 24'h0000ff;
		12'd1393: rd_data_0 <= 24'h0000ff;
		12'd1394: rd_data_0 <= 24'h0000ff;
		12'd1395: rd_data_0 <= 24'h0000ff;
		12'd1396: rd_data_0 <= 24'h0000ff;
		12'd1397: rd_data_0 <= 24'h0000ff;
		12'd1398: rd_data_0 <= 24'h0000ff;
		12'd1399: rd_data_0 <= 24'h0000ff;
		12'd1400: rd_data_0 <= 24'h000000;
		12'd1401: rd_data_0 <= 24'h000000;
		12'd1402: rd_data_0 <= 24'h000000;
		12'd1403: rd_data_0 <= 24'h000000;
		12'd1404: rd_data_0 <= 24'h000000;
		12'd1405: rd_data_0 <= 24'h000000;
		12'd1406: rd_data_0 <= 24'h000000;
		12'd1407: rd_data_0 <= 24'h000000;
		12'd1408: rd_data_0 <= 24'hffffff;
		12'd1409: rd_data_0 <= 24'hffffff;
		12'd1410: rd_data_0 <= 24'hffffff;
		12'd1411: rd_data_0 <= 24'hffffff;
		12'd1412: rd_data_0 <= 24'hffffff;
		12'd1413: rd_data_0 <= 24'hffffff;
		12'd1414: rd_data_0 <= 24'hffffff;
		12'd1415: rd_data_0 <= 24'hffffff;
		12'd1416: rd_data_0 <= 24'hffff00;
		12'd1417: rd_data_0 <= 24'hffff00;
		12'd1418: rd_data_0 <= 24'hffff00;
		12'd1419: rd_data_0 <= 24'hffff00;
		12'd1420: rd_data_0 <= 24'hffff00;
		12'd1421: rd_data_0 <= 24'hffff00;
		12'd1422: rd_data_0 <= 24'hffff00;
		12'd1423: rd_data_0 <= 24'hffff00;
		12'd1424: rd_data_0 <= 24'h00ffff;
		12'd1425: rd_data_0 <= 24'h00ffff;
		12'd1426: rd_data_0 <= 24'h00ffff;
		12'd1427: rd_data_0 <= 24'h00ffff;
		12'd1428: rd_data_0 <= 24'h00ffff;
		12'd1429: rd_data_0 <= 24'h00ffff;
		12'd1430: rd_data_0 <= 24'h00ffff;
		12'd1431: rd_data_0 <= 24'h00ffff;
		12'd1432: rd_data_0 <= 24'h00ff00;
		12'd1433: rd_data_0 <= 24'h00ff00;
		12'd1434: rd_data_0 <= 24'h00ff00;
		12'd1435: rd_data_0 <= 24'h00ff00;
		12'd1436: rd_data_0 <= 24'h00ff00;
		12'd1437: rd_data_0 <= 24'h00ff00;
		12'd1438: rd_data_0 <= 24'h00ff00;
		12'd1439: rd_data_0 <= 24'h00ff00;
		12'd1440: rd_data_0 <= 24'hff00ff;
		12'd1441: rd_data_0 <= 24'hff00ff;
		12'd1442: rd_data_0 <= 24'hff00ff;
		12'd1443: rd_data_0 <= 24'hff00ff;
		12'd1444: rd_data_0 <= 24'hff00ff;
		12'd1445: rd_data_0 <= 24'hff00ff;
		12'd1446: rd_data_0 <= 24'hff00ff;
		12'd1447: rd_data_0 <= 24'hff00ff;
		12'd1448: rd_data_0 <= 24'hff0000;
		12'd1449: rd_data_0 <= 24'hff0000;
		12'd1450: rd_data_0 <= 24'hff0000;
		12'd1451: rd_data_0 <= 24'hff0000;
		12'd1452: rd_data_0 <= 24'hff0000;
		12'd1453: rd_data_0 <= 24'hff0000;
		12'd1454: rd_data_0 <= 24'hff0000;
		12'd1455: rd_data_0 <= 24'hff0000;
		12'd1456: rd_data_0 <= 24'h0000ff;
		12'd1457: rd_data_0 <= 24'h0000ff;
		12'd1458: rd_data_0 <= 24'h0000ff;
		12'd1459: rd_data_0 <= 24'h0000ff;
		12'd1460: rd_data_0 <= 24'h0000ff;
		12'd1461: rd_data_0 <= 24'h0000ff;
		12'd1462: rd_data_0 <= 24'h0000ff;
		12'd1463: rd_data_0 <= 24'h0000ff;
		12'd1464: rd_data_0 <= 24'h000000;
		12'd1465: rd_data_0 <= 24'h000000;
		12'd1466: rd_data_0 <= 24'h000000;
		12'd1467: rd_data_0 <= 24'h000000;
		12'd1468: rd_data_0 <= 24'h000000;
		12'd1469: rd_data_0 <= 24'h000000;
		12'd1470: rd_data_0 <= 24'h000000;
		12'd1471: rd_data_0 <= 24'h000000;
		12'd1472: rd_data_0 <= 24'hffffff;
		12'd1473: rd_data_0 <= 24'hffffff;
		12'd1474: rd_data_0 <= 24'hffffff;
		12'd1475: rd_data_0 <= 24'hffffff;
		12'd1476: rd_data_0 <= 24'hffffff;
		12'd1477: rd_data_0 <= 24'hffffff;
		12'd1478: rd_data_0 <= 24'hffffff;
		12'd1479: rd_data_0 <= 24'hffffff;
		12'd1480: rd_data_0 <= 24'hffff00;
		12'd1481: rd_data_0 <= 24'hffff00;
		12'd1482: rd_data_0 <= 24'hffff00;
		12'd1483: rd_data_0 <= 24'hffff00;
		12'd1484: rd_data_0 <= 24'hffff00;
		12'd1485: rd_data_0 <= 24'hffff00;
		12'd1486: rd_data_0 <= 24'hffff00;
		12'd1487: rd_data_0 <= 24'hffff00;
		12'd1488: rd_data_0 <= 24'h00ffff;
		12'd1489: rd_data_0 <= 24'h00ffff;
		12'd1490: rd_data_0 <= 24'h00ffff;
		12'd1491: rd_data_0 <= 24'h00ffff;
		12'd1492: rd_data_0 <= 24'h00ffff;
		12'd1493: rd_data_0 <= 24'h00ffff;
		12'd1494: rd_data_0 <= 24'h00ffff;
		12'd1495: rd_data_0 <= 24'h00ffff;
		12'd1496: rd_data_0 <= 24'h00ff00;
		12'd1497: rd_data_0 <= 24'h00ff00;
		12'd1498: rd_data_0 <= 24'h00ff00;
		12'd1499: rd_data_0 <= 24'h00ff00;
		12'd1500: rd_data_0 <= 24'h00ff00;
		12'd1501: rd_data_0 <= 24'h00ff00;
		12'd1502: rd_data_0 <= 24'h00ff00;
		12'd1503: rd_data_0 <= 24'h00ff00;
		12'd1504: rd_data_0 <= 24'hff00ff;
		12'd1505: rd_data_0 <= 24'hff00ff;
		12'd1506: rd_data_0 <= 24'hff00ff;
		12'd1507: rd_data_0 <= 24'hff00ff;
		12'd1508: rd_data_0 <= 24'hff00ff;
		12'd1509: rd_data_0 <= 24'hff00ff;
		12'd1510: rd_data_0 <= 24'hff00ff;
		12'd1511: rd_data_0 <= 24'hff00ff;
		12'd1512: rd_data_0 <= 24'hff0000;
		12'd1513: rd_data_0 <= 24'hff0000;
		12'd1514: rd_data_0 <= 24'hff0000;
		12'd1515: rd_data_0 <= 24'hff0000;
		12'd1516: rd_data_0 <= 24'hff0000;
		12'd1517: rd_data_0 <= 24'hff0000;
		12'd1518: rd_data_0 <= 24'hff0000;
		12'd1519: rd_data_0 <= 24'hff0000;
		12'd1520: rd_data_0 <= 24'h0000ff;
		12'd1521: rd_data_0 <= 24'h0000ff;
		12'd1522: rd_data_0 <= 24'h0000ff;
		12'd1523: rd_data_0 <= 24'h0000ff;
		12'd1524: rd_data_0 <= 24'h0000ff;
		12'd1525: rd_data_0 <= 24'h0000ff;
		12'd1526: rd_data_0 <= 24'h0000ff;
		12'd1527: rd_data_0 <= 24'h0000ff;
		12'd1528: rd_data_0 <= 24'h000000;
		12'd1529: rd_data_0 <= 24'h000000;
		12'd1530: rd_data_0 <= 24'h000000;
		12'd1531: rd_data_0 <= 24'h000000;
		12'd1532: rd_data_0 <= 24'h000000;
		12'd1533: rd_data_0 <= 24'h000000;
		12'd1534: rd_data_0 <= 24'h000000;
		12'd1535: rd_data_0 <= 24'h000000;
		12'd1536: rd_data_0 <= 24'hffffff;
		12'd1537: rd_data_0 <= 24'hffffff;
		12'd1538: rd_data_0 <= 24'hffffff;
		12'd1539: rd_data_0 <= 24'hffffff;
		12'd1540: rd_data_0 <= 24'hffffff;
		12'd1541: rd_data_0 <= 24'hffffff;
		12'd1542: rd_data_0 <= 24'hffffff;
		12'd1543: rd_data_0 <= 24'hffffff;
		12'd1544: rd_data_0 <= 24'hffff00;
		12'd1545: rd_data_0 <= 24'hffff00;
		12'd1546: rd_data_0 <= 24'hffff00;
		12'd1547: rd_data_0 <= 24'hffff00;
		12'd1548: rd_data_0 <= 24'hffff00;
		12'd1549: rd_data_0 <= 24'hffff00;
		12'd1550: rd_data_0 <= 24'hffff00;
		12'd1551: rd_data_0 <= 24'hffff00;
		12'd1552: rd_data_0 <= 24'h00ffff;
		12'd1553: rd_data_0 <= 24'h00ffff;
		12'd1554: rd_data_0 <= 24'h00ffff;
		12'd1555: rd_data_0 <= 24'h00ffff;
		12'd1556: rd_data_0 <= 24'h00ffff;
		12'd1557: rd_data_0 <= 24'h00ffff;
		12'd1558: rd_data_0 <= 24'h00ffff;
		12'd1559: rd_data_0 <= 24'h00ffff;
		12'd1560: rd_data_0 <= 24'h00ff00;
		12'd1561: rd_data_0 <= 24'h00ff00;
		12'd1562: rd_data_0 <= 24'h00ff00;
		12'd1563: rd_data_0 <= 24'h00ff00;
		12'd1564: rd_data_0 <= 24'h00ff00;
		12'd1565: rd_data_0 <= 24'h00ff00;
		12'd1566: rd_data_0 <= 24'h00ff00;
		12'd1567: rd_data_0 <= 24'h00ff00;
		12'd1568: rd_data_0 <= 24'hff00ff;
		12'd1569: rd_data_0 <= 24'hff00ff;
		12'd1570: rd_data_0 <= 24'hff00ff;
		12'd1571: rd_data_0 <= 24'hff00ff;
		12'd1572: rd_data_0 <= 24'hff00ff;
		12'd1573: rd_data_0 <= 24'hff00ff;
		12'd1574: rd_data_0 <= 24'hff00ff;
		12'd1575: rd_data_0 <= 24'hff00ff;
		12'd1576: rd_data_0 <= 24'hff0000;
		12'd1577: rd_data_0 <= 24'hff0000;
		12'd1578: rd_data_0 <= 24'hff0000;
		12'd1579: rd_data_0 <= 24'hff0000;
		12'd1580: rd_data_0 <= 24'hff0000;
		12'd1581: rd_data_0 <= 24'hff0000;
		12'd1582: rd_data_0 <= 24'hff0000;
		12'd1583: rd_data_0 <= 24'hff0000;
		12'd1584: rd_data_0 <= 24'h0000ff;
		12'd1585: rd_data_0 <= 24'h0000ff;
		12'd1586: rd_data_0 <= 24'h0000ff;
		12'd1587: rd_data_0 <= 24'h0000ff;
		12'd1588: rd_data_0 <= 24'h0000ff;
		12'd1589: rd_data_0 <= 24'h0000ff;
		12'd1590: rd_data_0 <= 24'h0000ff;
		12'd1591: rd_data_0 <= 24'h0000ff;
		12'd1592: rd_data_0 <= 24'h000000;
		12'd1593: rd_data_0 <= 24'h000000;
		12'd1594: rd_data_0 <= 24'h000000;
		12'd1595: rd_data_0 <= 24'h000000;
		12'd1596: rd_data_0 <= 24'h000000;
		12'd1597: rd_data_0 <= 24'h000000;
		12'd1598: rd_data_0 <= 24'h000000;
		12'd1599: rd_data_0 <= 24'h000000;
		12'd1600: rd_data_0 <= 24'hffffff;
		12'd1601: rd_data_0 <= 24'hffffff;
		12'd1602: rd_data_0 <= 24'hffffff;
		12'd1603: rd_data_0 <= 24'hffffff;
		12'd1604: rd_data_0 <= 24'hffffff;
		12'd1605: rd_data_0 <= 24'hffffff;
		12'd1606: rd_data_0 <= 24'hffffff;
		12'd1607: rd_data_0 <= 24'hffffff;
		12'd1608: rd_data_0 <= 24'hffff00;
		12'd1609: rd_data_0 <= 24'hffff00;
		12'd1610: rd_data_0 <= 24'hffff00;
		12'd1611: rd_data_0 <= 24'hffff00;
		12'd1612: rd_data_0 <= 24'hffff00;
		12'd1613: rd_data_0 <= 24'hffff00;
		12'd1614: rd_data_0 <= 24'hffff00;
		12'd1615: rd_data_0 <= 24'hffff00;
		12'd1616: rd_data_0 <= 24'h00ffff;
		12'd1617: rd_data_0 <= 24'h00ffff;
		12'd1618: rd_data_0 <= 24'h00ffff;
		12'd1619: rd_data_0 <= 24'h00ffff;
		12'd1620: rd_data_0 <= 24'h00ffff;
		12'd1621: rd_data_0 <= 24'h00ffff;
		12'd1622: rd_data_0 <= 24'h00ffff;
		12'd1623: rd_data_0 <= 24'h00ffff;
		12'd1624: rd_data_0 <= 24'h00ff00;
		12'd1625: rd_data_0 <= 24'h00ff00;
		12'd1626: rd_data_0 <= 24'h00ff00;
		12'd1627: rd_data_0 <= 24'h00ff00;
		12'd1628: rd_data_0 <= 24'h00ff00;
		12'd1629: rd_data_0 <= 24'h00ff00;
		12'd1630: rd_data_0 <= 24'h00ff00;
		12'd1631: rd_data_0 <= 24'h00ff00;
		12'd1632: rd_data_0 <= 24'hff00ff;
		12'd1633: rd_data_0 <= 24'hff00ff;
		12'd1634: rd_data_0 <= 24'hff00ff;
		12'd1635: rd_data_0 <= 24'hff00ff;
		12'd1636: rd_data_0 <= 24'hff00ff;
		12'd1637: rd_data_0 <= 24'hff00ff;
		12'd1638: rd_data_0 <= 24'hff00ff;
		12'd1639: rd_data_0 <= 24'hff00ff;
		12'd1640: rd_data_0 <= 24'hff0000;
		12'd1641: rd_data_0 <= 24'hff0000;
		12'd1642: rd_data_0 <= 24'hff0000;
		12'd1643: rd_data_0 <= 24'hff0000;
		12'd1644: rd_data_0 <= 24'hff0000;
		12'd1645: rd_data_0 <= 24'hff0000;
		12'd1646: rd_data_0 <= 24'hff0000;
		12'd1647: rd_data_0 <= 24'hff0000;
		12'd1648: rd_data_0 <= 24'h0000ff;
		12'd1649: rd_data_0 <= 24'h0000ff;
		12'd1650: rd_data_0 <= 24'h0000ff;
		12'd1651: rd_data_0 <= 24'h0000ff;
		12'd1652: rd_data_0 <= 24'h0000ff;
		12'd1653: rd_data_0 <= 24'h0000ff;
		12'd1654: rd_data_0 <= 24'h0000ff;
		12'd1655: rd_data_0 <= 24'h0000ff;
		12'd1656: rd_data_0 <= 24'h000000;
		12'd1657: rd_data_0 <= 24'h000000;
		12'd1658: rd_data_0 <= 24'h000000;
		12'd1659: rd_data_0 <= 24'h000000;
		12'd1660: rd_data_0 <= 24'h000000;
		12'd1661: rd_data_0 <= 24'h000000;
		12'd1662: rd_data_0 <= 24'h000000;
		12'd1663: rd_data_0 <= 24'h000000;
		12'd1664: rd_data_0 <= 24'hffffff;
		12'd1665: rd_data_0 <= 24'hffffff;
		12'd1666: rd_data_0 <= 24'hffffff;
		12'd1667: rd_data_0 <= 24'hffffff;
		12'd1668: rd_data_0 <= 24'hffffff;
		12'd1669: rd_data_0 <= 24'hffffff;
		12'd1670: rd_data_0 <= 24'hffffff;
		12'd1671: rd_data_0 <= 24'hffffff;
		12'd1672: rd_data_0 <= 24'hffff00;
		12'd1673: rd_data_0 <= 24'hffff00;
		12'd1674: rd_data_0 <= 24'hffff00;
		12'd1675: rd_data_0 <= 24'hffff00;
		12'd1676: rd_data_0 <= 24'hffff00;
		12'd1677: rd_data_0 <= 24'hffff00;
		12'd1678: rd_data_0 <= 24'hffff00;
		12'd1679: rd_data_0 <= 24'hffff00;
		12'd1680: rd_data_0 <= 24'h00ffff;
		12'd1681: rd_data_0 <= 24'h00ffff;
		12'd1682: rd_data_0 <= 24'h00ffff;
		12'd1683: rd_data_0 <= 24'h00ffff;
		12'd1684: rd_data_0 <= 24'h00ffff;
		12'd1685: rd_data_0 <= 24'h00ffff;
		12'd1686: rd_data_0 <= 24'h00ffff;
		12'd1687: rd_data_0 <= 24'h00ffff;
		12'd1688: rd_data_0 <= 24'h00ff00;
		12'd1689: rd_data_0 <= 24'h00ff00;
		12'd1690: rd_data_0 <= 24'h00ff00;
		12'd1691: rd_data_0 <= 24'h00ff00;
		12'd1692: rd_data_0 <= 24'h00ff00;
		12'd1693: rd_data_0 <= 24'h00ff00;
		12'd1694: rd_data_0 <= 24'h00ff00;
		12'd1695: rd_data_0 <= 24'h00ff00;
		12'd1696: rd_data_0 <= 24'hff00ff;
		12'd1697: rd_data_0 <= 24'hff00ff;
		12'd1698: rd_data_0 <= 24'hff00ff;
		12'd1699: rd_data_0 <= 24'hff00ff;
		12'd1700: rd_data_0 <= 24'hff00ff;
		12'd1701: rd_data_0 <= 24'hff00ff;
		12'd1702: rd_data_0 <= 24'hff00ff;
		12'd1703: rd_data_0 <= 24'hff00ff;
		12'd1704: rd_data_0 <= 24'hff0000;
		12'd1705: rd_data_0 <= 24'hff0000;
		12'd1706: rd_data_0 <= 24'hff0000;
		12'd1707: rd_data_0 <= 24'hff0000;
		12'd1708: rd_data_0 <= 24'hff0000;
		12'd1709: rd_data_0 <= 24'hff0000;
		12'd1710: rd_data_0 <= 24'hff0000;
		12'd1711: rd_data_0 <= 24'hff0000;
		12'd1712: rd_data_0 <= 24'h0000ff;
		12'd1713: rd_data_0 <= 24'h0000ff;
		12'd1714: rd_data_0 <= 24'h0000ff;
		12'd1715: rd_data_0 <= 24'h0000ff;
		12'd1716: rd_data_0 <= 24'h0000ff;
		12'd1717: rd_data_0 <= 24'h0000ff;
		12'd1718: rd_data_0 <= 24'h0000ff;
		12'd1719: rd_data_0 <= 24'h0000ff;
		12'd1720: rd_data_0 <= 24'h000000;
		12'd1721: rd_data_0 <= 24'h000000;
		12'd1722: rd_data_0 <= 24'h000000;
		12'd1723: rd_data_0 <= 24'h000000;
		12'd1724: rd_data_0 <= 24'h000000;
		12'd1725: rd_data_0 <= 24'h000000;
		12'd1726: rd_data_0 <= 24'h000000;
		12'd1727: rd_data_0 <= 24'h000000;
		12'd1728: rd_data_0 <= 24'hffffff;
		12'd1729: rd_data_0 <= 24'hffffff;
		12'd1730: rd_data_0 <= 24'hffffff;
		12'd1731: rd_data_0 <= 24'hffffff;
		12'd1732: rd_data_0 <= 24'hffffff;
		12'd1733: rd_data_0 <= 24'hffffff;
		12'd1734: rd_data_0 <= 24'hffffff;
		12'd1735: rd_data_0 <= 24'hffffff;
		12'd1736: rd_data_0 <= 24'hffff00;
		12'd1737: rd_data_0 <= 24'hffff00;
		12'd1738: rd_data_0 <= 24'hffff00;
		12'd1739: rd_data_0 <= 24'hffff00;
		12'd1740: rd_data_0 <= 24'hffff00;
		12'd1741: rd_data_0 <= 24'hffff00;
		12'd1742: rd_data_0 <= 24'hffff00;
		12'd1743: rd_data_0 <= 24'hffff00;
		12'd1744: rd_data_0 <= 24'h00ffff;
		12'd1745: rd_data_0 <= 24'h00ffff;
		12'd1746: rd_data_0 <= 24'h00ffff;
		12'd1747: rd_data_0 <= 24'h00ffff;
		12'd1748: rd_data_0 <= 24'h00ffff;
		12'd1749: rd_data_0 <= 24'h00ffff;
		12'd1750: rd_data_0 <= 24'h00ffff;
		12'd1751: rd_data_0 <= 24'h00ffff;
		12'd1752: rd_data_0 <= 24'h00ff00;
		12'd1753: rd_data_0 <= 24'h00ff00;
		12'd1754: rd_data_0 <= 24'h00ff00;
		12'd1755: rd_data_0 <= 24'h00ff00;
		12'd1756: rd_data_0 <= 24'h00ff00;
		12'd1757: rd_data_0 <= 24'h00ff00;
		12'd1758: rd_data_0 <= 24'h00ff00;
		12'd1759: rd_data_0 <= 24'h00ff00;
		12'd1760: rd_data_0 <= 24'hff00ff;
		12'd1761: rd_data_0 <= 24'hff00ff;
		12'd1762: rd_data_0 <= 24'hff00ff;
		12'd1763: rd_data_0 <= 24'hff00ff;
		12'd1764: rd_data_0 <= 24'hff00ff;
		12'd1765: rd_data_0 <= 24'hff00ff;
		12'd1766: rd_data_0 <= 24'hff00ff;
		12'd1767: rd_data_0 <= 24'hff00ff;
		12'd1768: rd_data_0 <= 24'hff0000;
		12'd1769: rd_data_0 <= 24'hff0000;
		12'd1770: rd_data_0 <= 24'hff0000;
		12'd1771: rd_data_0 <= 24'hff0000;
		12'd1772: rd_data_0 <= 24'hff0000;
		12'd1773: rd_data_0 <= 24'hff0000;
		12'd1774: rd_data_0 <= 24'hff0000;
		12'd1775: rd_data_0 <= 24'hff0000;
		12'd1776: rd_data_0 <= 24'h0000ff;
		12'd1777: rd_data_0 <= 24'h0000ff;
		12'd1778: rd_data_0 <= 24'h0000ff;
		12'd1779: rd_data_0 <= 24'h0000ff;
		12'd1780: rd_data_0 <= 24'h0000ff;
		12'd1781: rd_data_0 <= 24'h0000ff;
		12'd1782: rd_data_0 <= 24'h0000ff;
		12'd1783: rd_data_0 <= 24'h0000ff;
		12'd1784: rd_data_0 <= 24'h000000;
		12'd1785: rd_data_0 <= 24'h000000;
		12'd1786: rd_data_0 <= 24'h000000;
		12'd1787: rd_data_0 <= 24'h000000;
		12'd1788: rd_data_0 <= 24'h000000;
		12'd1789: rd_data_0 <= 24'h000000;
		12'd1790: rd_data_0 <= 24'h000000;
		12'd1791: rd_data_0 <= 24'h000000;
		12'd1792: rd_data_0 <= 24'hffffff;
		12'd1793: rd_data_0 <= 24'hffffff;
		12'd1794: rd_data_0 <= 24'hffffff;
		12'd1795: rd_data_0 <= 24'hffffff;
		12'd1796: rd_data_0 <= 24'hffffff;
		12'd1797: rd_data_0 <= 24'hffffff;
		12'd1798: rd_data_0 <= 24'hffffff;
		12'd1799: rd_data_0 <= 24'hffffff;
		12'd1800: rd_data_0 <= 24'hffff00;
		12'd1801: rd_data_0 <= 24'hffff00;
		12'd1802: rd_data_0 <= 24'hffff00;
		12'd1803: rd_data_0 <= 24'hffff00;
		12'd1804: rd_data_0 <= 24'hffff00;
		12'd1805: rd_data_0 <= 24'hffff00;
		12'd1806: rd_data_0 <= 24'hffff00;
		12'd1807: rd_data_0 <= 24'hffff00;
		12'd1808: rd_data_0 <= 24'h00ffff;
		12'd1809: rd_data_0 <= 24'h00ffff;
		12'd1810: rd_data_0 <= 24'h00ffff;
		12'd1811: rd_data_0 <= 24'h00ffff;
		12'd1812: rd_data_0 <= 24'h00ffff;
		12'd1813: rd_data_0 <= 24'h00ffff;
		12'd1814: rd_data_0 <= 24'h00ffff;
		12'd1815: rd_data_0 <= 24'h00ffff;
		12'd1816: rd_data_0 <= 24'h00ff00;
		12'd1817: rd_data_0 <= 24'h00ff00;
		12'd1818: rd_data_0 <= 24'h00ff00;
		12'd1819: rd_data_0 <= 24'h00ff00;
		12'd1820: rd_data_0 <= 24'h00ff00;
		12'd1821: rd_data_0 <= 24'h00ff00;
		12'd1822: rd_data_0 <= 24'h00ff00;
		12'd1823: rd_data_0 <= 24'h00ff00;
		12'd1824: rd_data_0 <= 24'hff00ff;
		12'd1825: rd_data_0 <= 24'hff00ff;
		12'd1826: rd_data_0 <= 24'hff00ff;
		12'd1827: rd_data_0 <= 24'hff00ff;
		12'd1828: rd_data_0 <= 24'hff00ff;
		12'd1829: rd_data_0 <= 24'hff00ff;
		12'd1830: rd_data_0 <= 24'hff00ff;
		12'd1831: rd_data_0 <= 24'hff00ff;
		12'd1832: rd_data_0 <= 24'hff0000;
		12'd1833: rd_data_0 <= 24'hff0000;
		12'd1834: rd_data_0 <= 24'hff0000;
		12'd1835: rd_data_0 <= 24'hff0000;
		12'd1836: rd_data_0 <= 24'hff0000;
		12'd1837: rd_data_0 <= 24'hff0000;
		12'd1838: rd_data_0 <= 24'hff0000;
		12'd1839: rd_data_0 <= 24'hff0000;
		12'd1840: rd_data_0 <= 24'h0000ff;
		12'd1841: rd_data_0 <= 24'h0000ff;
		12'd1842: rd_data_0 <= 24'h0000ff;
		12'd1843: rd_data_0 <= 24'h0000ff;
		12'd1844: rd_data_0 <= 24'h0000ff;
		12'd1845: rd_data_0 <= 24'h0000ff;
		12'd1846: rd_data_0 <= 24'h0000ff;
		12'd1847: rd_data_0 <= 24'h0000ff;
		12'd1848: rd_data_0 <= 24'h000000;
		12'd1849: rd_data_0 <= 24'h000000;
		12'd1850: rd_data_0 <= 24'h000000;
		12'd1851: rd_data_0 <= 24'h000000;
		12'd1852: rd_data_0 <= 24'h000000;
		12'd1853: rd_data_0 <= 24'h000000;
		12'd1854: rd_data_0 <= 24'h000000;
		12'd1855: rd_data_0 <= 24'h000000;
		12'd1856: rd_data_0 <= 24'hffffff;
		12'd1857: rd_data_0 <= 24'hffffff;
		12'd1858: rd_data_0 <= 24'hffffff;
		12'd1859: rd_data_0 <= 24'hffffff;
		12'd1860: rd_data_0 <= 24'hffffff;
		12'd1861: rd_data_0 <= 24'hffffff;
		12'd1862: rd_data_0 <= 24'hffffff;
		12'd1863: rd_data_0 <= 24'hffffff;
		12'd1864: rd_data_0 <= 24'hffff00;
		12'd1865: rd_data_0 <= 24'hffff00;
		12'd1866: rd_data_0 <= 24'hffff00;
		12'd1867: rd_data_0 <= 24'hffff00;
		12'd1868: rd_data_0 <= 24'hffff00;
		12'd1869: rd_data_0 <= 24'hffff00;
		12'd1870: rd_data_0 <= 24'hffff00;
		12'd1871: rd_data_0 <= 24'hffff00;
		12'd1872: rd_data_0 <= 24'h00ffff;
		12'd1873: rd_data_0 <= 24'h00ffff;
		12'd1874: rd_data_0 <= 24'h00ffff;
		12'd1875: rd_data_0 <= 24'h00ffff;
		12'd1876: rd_data_0 <= 24'h00ffff;
		12'd1877: rd_data_0 <= 24'h00ffff;
		12'd1878: rd_data_0 <= 24'h00ffff;
		12'd1879: rd_data_0 <= 24'h00ffff;
		12'd1880: rd_data_0 <= 24'h00ff00;
		12'd1881: rd_data_0 <= 24'h00ff00;
		12'd1882: rd_data_0 <= 24'h00ff00;
		12'd1883: rd_data_0 <= 24'h00ff00;
		12'd1884: rd_data_0 <= 24'h00ff00;
		12'd1885: rd_data_0 <= 24'h00ff00;
		12'd1886: rd_data_0 <= 24'h00ff00;
		12'd1887: rd_data_0 <= 24'h00ff00;
		12'd1888: rd_data_0 <= 24'hff00ff;
		12'd1889: rd_data_0 <= 24'hff00ff;
		12'd1890: rd_data_0 <= 24'hff00ff;
		12'd1891: rd_data_0 <= 24'hff00ff;
		12'd1892: rd_data_0 <= 24'hff00ff;
		12'd1893: rd_data_0 <= 24'hff00ff;
		12'd1894: rd_data_0 <= 24'hff00ff;
		12'd1895: rd_data_0 <= 24'hff00ff;
		12'd1896: rd_data_0 <= 24'hff0000;
		12'd1897: rd_data_0 <= 24'hff0000;
		12'd1898: rd_data_0 <= 24'hff0000;
		12'd1899: rd_data_0 <= 24'hff0000;
		12'd1900: rd_data_0 <= 24'hff0000;
		12'd1901: rd_data_0 <= 24'hff0000;
		12'd1902: rd_data_0 <= 24'hff0000;
		12'd1903: rd_data_0 <= 24'hff0000;
		12'd1904: rd_data_0 <= 24'h0000ff;
		12'd1905: rd_data_0 <= 24'h0000ff;
		12'd1906: rd_data_0 <= 24'h0000ff;
		12'd1907: rd_data_0 <= 24'h0000ff;
		12'd1908: rd_data_0 <= 24'h0000ff;
		12'd1909: rd_data_0 <= 24'h0000ff;
		12'd1910: rd_data_0 <= 24'h0000ff;
		12'd1911: rd_data_0 <= 24'h0000ff;
		12'd1912: rd_data_0 <= 24'h000000;
		12'd1913: rd_data_0 <= 24'h000000;
		12'd1914: rd_data_0 <= 24'h000000;
		12'd1915: rd_data_0 <= 24'h000000;
		12'd1916: rd_data_0 <= 24'h000000;
		12'd1917: rd_data_0 <= 24'h000000;
		12'd1918: rd_data_0 <= 24'h000000;
		12'd1919: rd_data_0 <= 24'h000000;
		12'd1920: rd_data_0 <= 24'hffffff;
		12'd1921: rd_data_0 <= 24'hffffff;
		12'd1922: rd_data_0 <= 24'hffffff;
		12'd1923: rd_data_0 <= 24'hffffff;
		12'd1924: rd_data_0 <= 24'hffffff;
		12'd1925: rd_data_0 <= 24'hffffff;
		12'd1926: rd_data_0 <= 24'hffffff;
		12'd1927: rd_data_0 <= 24'hffffff;
		12'd1928: rd_data_0 <= 24'hffff00;
		12'd1929: rd_data_0 <= 24'hffff00;
		12'd1930: rd_data_0 <= 24'hffff00;
		12'd1931: rd_data_0 <= 24'hffff00;
		12'd1932: rd_data_0 <= 24'hffff00;
		12'd1933: rd_data_0 <= 24'hffff00;
		12'd1934: rd_data_0 <= 24'hffff00;
		12'd1935: rd_data_0 <= 24'hffff00;
		12'd1936: rd_data_0 <= 24'h00ffff;
		12'd1937: rd_data_0 <= 24'h00ffff;
		12'd1938: rd_data_0 <= 24'h00ffff;
		12'd1939: rd_data_0 <= 24'h00ffff;
		12'd1940: rd_data_0 <= 24'h00ffff;
		12'd1941: rd_data_0 <= 24'h00ffff;
		12'd1942: rd_data_0 <= 24'h00ffff;
		12'd1943: rd_data_0 <= 24'h00ffff;
		12'd1944: rd_data_0 <= 24'h00ff00;
		12'd1945: rd_data_0 <= 24'h00ff00;
		12'd1946: rd_data_0 <= 24'h00ff00;
		12'd1947: rd_data_0 <= 24'h00ff00;
		12'd1948: rd_data_0 <= 24'h00ff00;
		12'd1949: rd_data_0 <= 24'h00ff00;
		12'd1950: rd_data_0 <= 24'h00ff00;
		12'd1951: rd_data_0 <= 24'h00ff00;
		12'd1952: rd_data_0 <= 24'hff00ff;
		12'd1953: rd_data_0 <= 24'hff00ff;
		12'd1954: rd_data_0 <= 24'hff00ff;
		12'd1955: rd_data_0 <= 24'hff00ff;
		12'd1956: rd_data_0 <= 24'hff00ff;
		12'd1957: rd_data_0 <= 24'hff00ff;
		12'd1958: rd_data_0 <= 24'hff00ff;
		12'd1959: rd_data_0 <= 24'hff00ff;
		12'd1960: rd_data_0 <= 24'hff0000;
		12'd1961: rd_data_0 <= 24'hff0000;
		12'd1962: rd_data_0 <= 24'hff0000;
		12'd1963: rd_data_0 <= 24'hff0000;
		12'd1964: rd_data_0 <= 24'hff0000;
		12'd1965: rd_data_0 <= 24'hff0000;
		12'd1966: rd_data_0 <= 24'hff0000;
		12'd1967: rd_data_0 <= 24'hff0000;
		12'd1968: rd_data_0 <= 24'h0000ff;
		12'd1969: rd_data_0 <= 24'h0000ff;
		12'd1970: rd_data_0 <= 24'h0000ff;
		12'd1971: rd_data_0 <= 24'h0000ff;
		12'd1972: rd_data_0 <= 24'h0000ff;
		12'd1973: rd_data_0 <= 24'h0000ff;
		12'd1974: rd_data_0 <= 24'h0000ff;
		12'd1975: rd_data_0 <= 24'h0000ff;
		12'd1976: rd_data_0 <= 24'h000000;
		12'd1977: rd_data_0 <= 24'h000000;
		12'd1978: rd_data_0 <= 24'h000000;
		12'd1979: rd_data_0 <= 24'h000000;
		12'd1980: rd_data_0 <= 24'h000000;
		12'd1981: rd_data_0 <= 24'h000000;
		12'd1982: rd_data_0 <= 24'h000000;
		12'd1983: rd_data_0 <= 24'h000000;
		12'd1984: rd_data_0 <= 24'hffffff;
		12'd1985: rd_data_0 <= 24'hffffff;
		12'd1986: rd_data_0 <= 24'hffffff;
		12'd1987: rd_data_0 <= 24'hffffff;
		12'd1988: rd_data_0 <= 24'hffffff;
		12'd1989: rd_data_0 <= 24'hffffff;
		12'd1990: rd_data_0 <= 24'hffffff;
		12'd1991: rd_data_0 <= 24'hffffff;
		12'd1992: rd_data_0 <= 24'hffff00;
		12'd1993: rd_data_0 <= 24'hffff00;
		12'd1994: rd_data_0 <= 24'hffff00;
		12'd1995: rd_data_0 <= 24'hffff00;
		12'd1996: rd_data_0 <= 24'hffff00;
		12'd1997: rd_data_0 <= 24'hffff00;
		12'd1998: rd_data_0 <= 24'hffff00;
		12'd1999: rd_data_0 <= 24'hffff00;
		12'd2000: rd_data_0 <= 24'h00ffff;
		12'd2001: rd_data_0 <= 24'h00ffff;
		12'd2002: rd_data_0 <= 24'h00ffff;
		12'd2003: rd_data_0 <= 24'h00ffff;
		12'd2004: rd_data_0 <= 24'h00ffff;
		12'd2005: rd_data_0 <= 24'h00ffff;
		12'd2006: rd_data_0 <= 24'h00ffff;
		12'd2007: rd_data_0 <= 24'h00ffff;
		12'd2008: rd_data_0 <= 24'h00ff00;
		12'd2009: rd_data_0 <= 24'h00ff00;
		12'd2010: rd_data_0 <= 24'h00ff00;
		12'd2011: rd_data_0 <= 24'h00ff00;
		12'd2012: rd_data_0 <= 24'h00ff00;
		12'd2013: rd_data_0 <= 24'h00ff00;
		12'd2014: rd_data_0 <= 24'h00ff00;
		12'd2015: rd_data_0 <= 24'h00ff00;
		12'd2016: rd_data_0 <= 24'hff00ff;
		12'd2017: rd_data_0 <= 24'hff00ff;
		12'd2018: rd_data_0 <= 24'hff00ff;
		12'd2019: rd_data_0 <= 24'hff00ff;
		12'd2020: rd_data_0 <= 24'hff00ff;
		12'd2021: rd_data_0 <= 24'hff00ff;
		12'd2022: rd_data_0 <= 24'hff00ff;
		12'd2023: rd_data_0 <= 24'hff00ff;
		12'd2024: rd_data_0 <= 24'hff0000;
		12'd2025: rd_data_0 <= 24'hff0000;
		12'd2026: rd_data_0 <= 24'hff0000;
		12'd2027: rd_data_0 <= 24'hff0000;
		12'd2028: rd_data_0 <= 24'hff0000;
		12'd2029: rd_data_0 <= 24'hff0000;
		12'd2030: rd_data_0 <= 24'hff0000;
		12'd2031: rd_data_0 <= 24'hff0000;
		12'd2032: rd_data_0 <= 24'h0000ff;
		12'd2033: rd_data_0 <= 24'h0000ff;
		12'd2034: rd_data_0 <= 24'h0000ff;
		12'd2035: rd_data_0 <= 24'h0000ff;
		12'd2036: rd_data_0 <= 24'h0000ff;
		12'd2037: rd_data_0 <= 24'h0000ff;
		12'd2038: rd_data_0 <= 24'h0000ff;
		12'd2039: rd_data_0 <= 24'h0000ff;
		12'd2040: rd_data_0 <= 24'h000000;
		12'd2041: rd_data_0 <= 24'h000000;
		12'd2042: rd_data_0 <= 24'h000000;
		12'd2043: rd_data_0 <= 24'h000000;
		12'd2044: rd_data_0 <= 24'h000000;
		12'd2045: rd_data_0 <= 24'h000000;
		12'd2046: rd_data_0 <= 24'h000000;
		12'd2047: rd_data_0 <= 24'h000000;

        endcase

        case (i_rd_addr)
		12'd0000: rd_data_1 <= 24'hffffff;
		12'd0001: rd_data_1 <= 24'hffffff;
		12'd0002: rd_data_1 <= 24'hffffff;
		12'd0003: rd_data_1 <= 24'hffffff;
		12'd0004: rd_data_1 <= 24'hffffff;
		12'd0005: rd_data_1 <= 24'hffffff;
		12'd0006: rd_data_1 <= 24'hffffff;
		12'd0007: rd_data_1 <= 24'hffffff;
		12'd0008: rd_data_1 <= 24'hffff00;
		12'd0009: rd_data_1 <= 24'hffff00;
		12'd0010: rd_data_1 <= 24'hffff00;
		12'd0011: rd_data_1 <= 24'hffff00;
		12'd0012: rd_data_1 <= 24'hffff00;
		12'd0013: rd_data_1 <= 24'hffff00;
		12'd0014: rd_data_1 <= 24'hffff00;
		12'd0015: rd_data_1 <= 24'hffff00;
		12'd0016: rd_data_1 <= 24'h00ffff;
		12'd0017: rd_data_1 <= 24'h00ffff;
		12'd0018: rd_data_1 <= 24'h00ffff;
		12'd0019: rd_data_1 <= 24'h00ffff;
		12'd0020: rd_data_1 <= 24'h00ffff;
		12'd0021: rd_data_1 <= 24'h00ffff;
		12'd0022: rd_data_1 <= 24'h00ffff;
		12'd0023: rd_data_1 <= 24'h00ffff;
		12'd0024: rd_data_1 <= 24'h00ff00;
		12'd0025: rd_data_1 <= 24'h00ff00;
		12'd0026: rd_data_1 <= 24'h00ff00;
		12'd0027: rd_data_1 <= 24'h00ff00;
		12'd0028: rd_data_1 <= 24'h00ff00;
		12'd0029: rd_data_1 <= 24'h00ff00;
		12'd0030: rd_data_1 <= 24'h00ff00;
		12'd0031: rd_data_1 <= 24'h00ff00;
		12'd0032: rd_data_1 <= 24'hff00ff;
		12'd0033: rd_data_1 <= 24'hff00ff;
		12'd0034: rd_data_1 <= 24'hff00ff;
		12'd0035: rd_data_1 <= 24'hff00ff;
		12'd0036: rd_data_1 <= 24'hff00ff;
		12'd0037: rd_data_1 <= 24'hff00ff;
		12'd0038: rd_data_1 <= 24'hff00ff;
		12'd0039: rd_data_1 <= 24'hff00ff;
		12'd0040: rd_data_1 <= 24'hff0000;
		12'd0041: rd_data_1 <= 24'hff0000;
		12'd0042: rd_data_1 <= 24'hff0000;
		12'd0043: rd_data_1 <= 24'hff0000;
		12'd0044: rd_data_1 <= 24'hff0000;
		12'd0045: rd_data_1 <= 24'hff0000;
		12'd0046: rd_data_1 <= 24'hff0000;
		12'd0047: rd_data_1 <= 24'hff0000;
		12'd0048: rd_data_1 <= 24'h0000ff;
		12'd0049: rd_data_1 <= 24'h0000ff;
		12'd0050: rd_data_1 <= 24'h0000ff;
		12'd0051: rd_data_1 <= 24'h0000ff;
		12'd0052: rd_data_1 <= 24'h0000ff;
		12'd0053: rd_data_1 <= 24'h0000ff;
		12'd0054: rd_data_1 <= 24'h0000ff;
		12'd0055: rd_data_1 <= 24'h0000ff;
		12'd0056: rd_data_1 <= 24'h000000;
		12'd0057: rd_data_1 <= 24'h000000;
		12'd0058: rd_data_1 <= 24'h000000;
		12'd0059: rd_data_1 <= 24'h000000;
		12'd0060: rd_data_1 <= 24'h000000;
		12'd0061: rd_data_1 <= 24'h000000;
		12'd0062: rd_data_1 <= 24'h000000;
		12'd0063: rd_data_1 <= 24'h000000;
		12'd0064: rd_data_1 <= 24'hffffff;
		12'd0065: rd_data_1 <= 24'hffffff;
		12'd0066: rd_data_1 <= 24'hffffff;
		12'd0067: rd_data_1 <= 24'hffffff;
		12'd0068: rd_data_1 <= 24'hffffff;
		12'd0069: rd_data_1 <= 24'hffffff;
		12'd0070: rd_data_1 <= 24'hffffff;
		12'd0071: rd_data_1 <= 24'hffffff;
		12'd0072: rd_data_1 <= 24'hffff00;
		12'd0073: rd_data_1 <= 24'hffff00;
		12'd0074: rd_data_1 <= 24'hffff00;
		12'd0075: rd_data_1 <= 24'hffff00;
		12'd0076: rd_data_1 <= 24'hffff00;
		12'd0077: rd_data_1 <= 24'hffff00;
		12'd0078: rd_data_1 <= 24'hffff00;
		12'd0079: rd_data_1 <= 24'hffff00;
		12'd0080: rd_data_1 <= 24'h00ffff;
		12'd0081: rd_data_1 <= 24'h00ffff;
		12'd0082: rd_data_1 <= 24'h00ffff;
		12'd0083: rd_data_1 <= 24'h00ffff;
		12'd0084: rd_data_1 <= 24'h00ffff;
		12'd0085: rd_data_1 <= 24'h00ffff;
		12'd0086: rd_data_1 <= 24'h00ffff;
		12'd0087: rd_data_1 <= 24'h00ffff;
		12'd0088: rd_data_1 <= 24'h00ff00;
		12'd0089: rd_data_1 <= 24'h00ff00;
		12'd0090: rd_data_1 <= 24'h00ff00;
		12'd0091: rd_data_1 <= 24'h00ff00;
		12'd0092: rd_data_1 <= 24'h00ff00;
		12'd0093: rd_data_1 <= 24'h00ff00;
		12'd0094: rd_data_1 <= 24'h00ff00;
		12'd0095: rd_data_1 <= 24'h00ff00;
		12'd0096: rd_data_1 <= 24'hff00ff;
		12'd0097: rd_data_1 <= 24'hff00ff;
		12'd0098: rd_data_1 <= 24'hff00ff;
		12'd0099: rd_data_1 <= 24'hff00ff;
		12'd0100: rd_data_1 <= 24'hff00ff;
		12'd0101: rd_data_1 <= 24'hff00ff;
		12'd0102: rd_data_1 <= 24'hff00ff;
		12'd0103: rd_data_1 <= 24'hff00ff;
		12'd0104: rd_data_1 <= 24'hff0000;
		12'd0105: rd_data_1 <= 24'hff0000;
		12'd0106: rd_data_1 <= 24'hff0000;
		12'd0107: rd_data_1 <= 24'hff0000;
		12'd0108: rd_data_1 <= 24'hff0000;
		12'd0109: rd_data_1 <= 24'hff0000;
		12'd0110: rd_data_1 <= 24'hff0000;
		12'd0111: rd_data_1 <= 24'hff0000;
		12'd0112: rd_data_1 <= 24'h0000ff;
		12'd0113: rd_data_1 <= 24'h0000ff;
		12'd0114: rd_data_1 <= 24'h0000ff;
		12'd0115: rd_data_1 <= 24'h0000ff;
		12'd0116: rd_data_1 <= 24'h0000ff;
		12'd0117: rd_data_1 <= 24'h0000ff;
		12'd0118: rd_data_1 <= 24'h0000ff;
		12'd0119: rd_data_1 <= 24'h0000ff;
		12'd0120: rd_data_1 <= 24'h000000;
		12'd0121: rd_data_1 <= 24'h000000;
		12'd0122: rd_data_1 <= 24'h000000;
		12'd0123: rd_data_1 <= 24'h000000;
		12'd0124: rd_data_1 <= 24'h000000;
		12'd0125: rd_data_1 <= 24'h000000;
		12'd0126: rd_data_1 <= 24'h000000;
		12'd0127: rd_data_1 <= 24'h000000;
		12'd0128: rd_data_1 <= 24'hffffff;
		12'd0129: rd_data_1 <= 24'hffffff;
		12'd0130: rd_data_1 <= 24'hffffff;
		12'd0131: rd_data_1 <= 24'hffffff;
		12'd0132: rd_data_1 <= 24'hffffff;
		12'd0133: rd_data_1 <= 24'hffffff;
		12'd0134: rd_data_1 <= 24'hffffff;
		12'd0135: rd_data_1 <= 24'hffffff;
		12'd0136: rd_data_1 <= 24'hffff00;
		12'd0137: rd_data_1 <= 24'hffff00;
		12'd0138: rd_data_1 <= 24'hffff00;
		12'd0139: rd_data_1 <= 24'hffff00;
		12'd0140: rd_data_1 <= 24'hffff00;
		12'd0141: rd_data_1 <= 24'hffff00;
		12'd0142: rd_data_1 <= 24'hffff00;
		12'd0143: rd_data_1 <= 24'hffff00;
		12'd0144: rd_data_1 <= 24'h00ffff;
		12'd0145: rd_data_1 <= 24'h00ffff;
		12'd0146: rd_data_1 <= 24'h00ffff;
		12'd0147: rd_data_1 <= 24'h00ffff;
		12'd0148: rd_data_1 <= 24'h00ffff;
		12'd0149: rd_data_1 <= 24'h00ffff;
		12'd0150: rd_data_1 <= 24'h00ffff;
		12'd0151: rd_data_1 <= 24'h00ffff;
		12'd0152: rd_data_1 <= 24'h00ff00;
		12'd0153: rd_data_1 <= 24'h00ff00;
		12'd0154: rd_data_1 <= 24'h00ff00;
		12'd0155: rd_data_1 <= 24'h00ff00;
		12'd0156: rd_data_1 <= 24'h00ff00;
		12'd0157: rd_data_1 <= 24'h00ff00;
		12'd0158: rd_data_1 <= 24'h00ff00;
		12'd0159: rd_data_1 <= 24'h00ff00;
		12'd0160: rd_data_1 <= 24'hff00ff;
		12'd0161: rd_data_1 <= 24'hff00ff;
		12'd0162: rd_data_1 <= 24'hff00ff;
		12'd0163: rd_data_1 <= 24'hff00ff;
		12'd0164: rd_data_1 <= 24'hff00ff;
		12'd0165: rd_data_1 <= 24'hff00ff;
		12'd0166: rd_data_1 <= 24'hff00ff;
		12'd0167: rd_data_1 <= 24'hff00ff;
		12'd0168: rd_data_1 <= 24'hff0000;
		12'd0169: rd_data_1 <= 24'hff0000;
		12'd0170: rd_data_1 <= 24'hff0000;
		12'd0171: rd_data_1 <= 24'hff0000;
		12'd0172: rd_data_1 <= 24'hff0000;
		12'd0173: rd_data_1 <= 24'hff0000;
		12'd0174: rd_data_1 <= 24'hff0000;
		12'd0175: rd_data_1 <= 24'hff0000;
		12'd0176: rd_data_1 <= 24'h0000ff;
		12'd0177: rd_data_1 <= 24'h0000ff;
		12'd0178: rd_data_1 <= 24'h0000ff;
		12'd0179: rd_data_1 <= 24'h0000ff;
		12'd0180: rd_data_1 <= 24'h0000ff;
		12'd0181: rd_data_1 <= 24'h0000ff;
		12'd0182: rd_data_1 <= 24'h0000ff;
		12'd0183: rd_data_1 <= 24'h0000ff;
		12'd0184: rd_data_1 <= 24'h000000;
		12'd0185: rd_data_1 <= 24'h000000;
		12'd0186: rd_data_1 <= 24'h000000;
		12'd0187: rd_data_1 <= 24'h000000;
		12'd0188: rd_data_1 <= 24'h000000;
		12'd0189: rd_data_1 <= 24'h000000;
		12'd0190: rd_data_1 <= 24'h000000;
		12'd0191: rd_data_1 <= 24'h000000;
		12'd0192: rd_data_1 <= 24'hffffff;
		12'd0193: rd_data_1 <= 24'hffffff;
		12'd0194: rd_data_1 <= 24'hffffff;
		12'd0195: rd_data_1 <= 24'hffffff;
		12'd0196: rd_data_1 <= 24'hffffff;
		12'd0197: rd_data_1 <= 24'hffffff;
		12'd0198: rd_data_1 <= 24'hffffff;
		12'd0199: rd_data_1 <= 24'hffffff;
		12'd0200: rd_data_1 <= 24'hffff00;
		12'd0201: rd_data_1 <= 24'hffff00;
		12'd0202: rd_data_1 <= 24'hffff00;
		12'd0203: rd_data_1 <= 24'hffff00;
		12'd0204: rd_data_1 <= 24'hffff00;
		12'd0205: rd_data_1 <= 24'hffff00;
		12'd0206: rd_data_1 <= 24'hffff00;
		12'd0207: rd_data_1 <= 24'hffff00;
		12'd0208: rd_data_1 <= 24'h00ffff;
		12'd0209: rd_data_1 <= 24'h00ffff;
		12'd0210: rd_data_1 <= 24'h00ffff;
		12'd0211: rd_data_1 <= 24'h00ffff;
		12'd0212: rd_data_1 <= 24'h00ffff;
		12'd0213: rd_data_1 <= 24'h00ffff;
		12'd0214: rd_data_1 <= 24'h00ffff;
		12'd0215: rd_data_1 <= 24'h00ffff;
		12'd0216: rd_data_1 <= 24'h00ff00;
		12'd0217: rd_data_1 <= 24'h00ff00;
		12'd0218: rd_data_1 <= 24'h00ff00;
		12'd0219: rd_data_1 <= 24'h00ff00;
		12'd0220: rd_data_1 <= 24'h00ff00;
		12'd0221: rd_data_1 <= 24'h00ff00;
		12'd0222: rd_data_1 <= 24'h00ff00;
		12'd0223: rd_data_1 <= 24'h00ff00;
		12'd0224: rd_data_1 <= 24'hff00ff;
		12'd0225: rd_data_1 <= 24'hff00ff;
		12'd0226: rd_data_1 <= 24'hff00ff;
		12'd0227: rd_data_1 <= 24'hff00ff;
		12'd0228: rd_data_1 <= 24'hff00ff;
		12'd0229: rd_data_1 <= 24'hff00ff;
		12'd0230: rd_data_1 <= 24'hff00ff;
		12'd0231: rd_data_1 <= 24'hff00ff;
		12'd0232: rd_data_1 <= 24'hff0000;
		12'd0233: rd_data_1 <= 24'hff0000;
		12'd0234: rd_data_1 <= 24'hff0000;
		12'd0235: rd_data_1 <= 24'hff0000;
		12'd0236: rd_data_1 <= 24'hff0000;
		12'd0237: rd_data_1 <= 24'hff0000;
		12'd0238: rd_data_1 <= 24'hff0000;
		12'd0239: rd_data_1 <= 24'hff0000;
		12'd0240: rd_data_1 <= 24'h0000ff;
		12'd0241: rd_data_1 <= 24'h0000ff;
		12'd0242: rd_data_1 <= 24'h0000ff;
		12'd0243: rd_data_1 <= 24'h0000ff;
		12'd0244: rd_data_1 <= 24'h0000ff;
		12'd0245: rd_data_1 <= 24'h0000ff;
		12'd0246: rd_data_1 <= 24'h0000ff;
		12'd0247: rd_data_1 <= 24'h0000ff;
		12'd0248: rd_data_1 <= 24'h000000;
		12'd0249: rd_data_1 <= 24'h000000;
		12'd0250: rd_data_1 <= 24'h000000;
		12'd0251: rd_data_1 <= 24'h000000;
		12'd0252: rd_data_1 <= 24'h000000;
		12'd0253: rd_data_1 <= 24'h000000;
		12'd0254: rd_data_1 <= 24'h000000;
		12'd0255: rd_data_1 <= 24'h000000;
		12'd0256: rd_data_1 <= 24'hffffff;
		12'd0257: rd_data_1 <= 24'hffffff;
		12'd0258: rd_data_1 <= 24'hffffff;
		12'd0259: rd_data_1 <= 24'hffffff;
		12'd0260: rd_data_1 <= 24'hffffff;
		12'd0261: rd_data_1 <= 24'hffffff;
		12'd0262: rd_data_1 <= 24'hffffff;
		12'd0263: rd_data_1 <= 24'hffffff;
		12'd0264: rd_data_1 <= 24'hffff00;
		12'd0265: rd_data_1 <= 24'hffff00;
		12'd0266: rd_data_1 <= 24'hffff00;
		12'd0267: rd_data_1 <= 24'hffff00;
		12'd0268: rd_data_1 <= 24'hffff00;
		12'd0269: rd_data_1 <= 24'hffff00;
		12'd0270: rd_data_1 <= 24'hffff00;
		12'd0271: rd_data_1 <= 24'hffff00;
		12'd0272: rd_data_1 <= 24'h00ffff;
		12'd0273: rd_data_1 <= 24'h00ffff;
		12'd0274: rd_data_1 <= 24'h00ffff;
		12'd0275: rd_data_1 <= 24'h00ffff;
		12'd0276: rd_data_1 <= 24'h00ffff;
		12'd0277: rd_data_1 <= 24'h00ffff;
		12'd0278: rd_data_1 <= 24'h00ffff;
		12'd0279: rd_data_1 <= 24'h00ffff;
		12'd0280: rd_data_1 <= 24'h00ff00;
		12'd0281: rd_data_1 <= 24'h00ff00;
		12'd0282: rd_data_1 <= 24'h00ff00;
		12'd0283: rd_data_1 <= 24'h00ff00;
		12'd0284: rd_data_1 <= 24'h00ff00;
		12'd0285: rd_data_1 <= 24'h00ff00;
		12'd0286: rd_data_1 <= 24'h00ff00;
		12'd0287: rd_data_1 <= 24'h00ff00;
		12'd0288: rd_data_1 <= 24'hff00ff;
		12'd0289: rd_data_1 <= 24'hff00ff;
		12'd0290: rd_data_1 <= 24'hff00ff;
		12'd0291: rd_data_1 <= 24'hff00ff;
		12'd0292: rd_data_1 <= 24'hff00ff;
		12'd0293: rd_data_1 <= 24'hff00ff;
		12'd0294: rd_data_1 <= 24'hff00ff;
		12'd0295: rd_data_1 <= 24'hff00ff;
		12'd0296: rd_data_1 <= 24'hff0000;
		12'd0297: rd_data_1 <= 24'hff0000;
		12'd0298: rd_data_1 <= 24'hff0000;
		12'd0299: rd_data_1 <= 24'hff0000;
		12'd0300: rd_data_1 <= 24'hff0000;
		12'd0301: rd_data_1 <= 24'hff0000;
		12'd0302: rd_data_1 <= 24'hff0000;
		12'd0303: rd_data_1 <= 24'hff0000;
		12'd0304: rd_data_1 <= 24'h0000ff;
		12'd0305: rd_data_1 <= 24'h0000ff;
		12'd0306: rd_data_1 <= 24'h0000ff;
		12'd0307: rd_data_1 <= 24'h0000ff;
		12'd0308: rd_data_1 <= 24'h0000ff;
		12'd0309: rd_data_1 <= 24'h0000ff;
		12'd0310: rd_data_1 <= 24'h0000ff;
		12'd0311: rd_data_1 <= 24'h0000ff;
		12'd0312: rd_data_1 <= 24'h000000;
		12'd0313: rd_data_1 <= 24'h000000;
		12'd0314: rd_data_1 <= 24'h000000;
		12'd0315: rd_data_1 <= 24'h000000;
		12'd0316: rd_data_1 <= 24'h000000;
		12'd0317: rd_data_1 <= 24'h000000;
		12'd0318: rd_data_1 <= 24'h000000;
		12'd0319: rd_data_1 <= 24'h000000;
		12'd0320: rd_data_1 <= 24'hffffff;
		12'd0321: rd_data_1 <= 24'hffffff;
		12'd0322: rd_data_1 <= 24'hffffff;
		12'd0323: rd_data_1 <= 24'hffffff;
		12'd0324: rd_data_1 <= 24'hffffff;
		12'd0325: rd_data_1 <= 24'hffffff;
		12'd0326: rd_data_1 <= 24'hffffff;
		12'd0327: rd_data_1 <= 24'hffffff;
		12'd0328: rd_data_1 <= 24'hffff00;
		12'd0329: rd_data_1 <= 24'hffff00;
		12'd0330: rd_data_1 <= 24'hffff00;
		12'd0331: rd_data_1 <= 24'hffff00;
		12'd0332: rd_data_1 <= 24'hffff00;
		12'd0333: rd_data_1 <= 24'hffff00;
		12'd0334: rd_data_1 <= 24'hffff00;
		12'd0335: rd_data_1 <= 24'hffff00;
		12'd0336: rd_data_1 <= 24'h00ffff;
		12'd0337: rd_data_1 <= 24'h00ffff;
		12'd0338: rd_data_1 <= 24'h00ffff;
		12'd0339: rd_data_1 <= 24'h00ffff;
		12'd0340: rd_data_1 <= 24'h00ffff;
		12'd0341: rd_data_1 <= 24'h00ffff;
		12'd0342: rd_data_1 <= 24'h00ffff;
		12'd0343: rd_data_1 <= 24'h00ffff;
		12'd0344: rd_data_1 <= 24'h00ff00;
		12'd0345: rd_data_1 <= 24'h00ff00;
		12'd0346: rd_data_1 <= 24'h00ff00;
		12'd0347: rd_data_1 <= 24'h00ff00;
		12'd0348: rd_data_1 <= 24'h00ff00;
		12'd0349: rd_data_1 <= 24'h00ff00;
		12'd0350: rd_data_1 <= 24'h00ff00;
		12'd0351: rd_data_1 <= 24'h00ff00;
		12'd0352: rd_data_1 <= 24'hff00ff;
		12'd0353: rd_data_1 <= 24'hff00ff;
		12'd0354: rd_data_1 <= 24'hff00ff;
		12'd0355: rd_data_1 <= 24'hff00ff;
		12'd0356: rd_data_1 <= 24'hff00ff;
		12'd0357: rd_data_1 <= 24'hff00ff;
		12'd0358: rd_data_1 <= 24'hff00ff;
		12'd0359: rd_data_1 <= 24'hff00ff;
		12'd0360: rd_data_1 <= 24'hff0000;
		12'd0361: rd_data_1 <= 24'hff0000;
		12'd0362: rd_data_1 <= 24'hff0000;
		12'd0363: rd_data_1 <= 24'hff0000;
		12'd0364: rd_data_1 <= 24'hff0000;
		12'd0365: rd_data_1 <= 24'hff0000;
		12'd0366: rd_data_1 <= 24'hff0000;
		12'd0367: rd_data_1 <= 24'hff0000;
		12'd0368: rd_data_1 <= 24'h0000ff;
		12'd0369: rd_data_1 <= 24'h0000ff;
		12'd0370: rd_data_1 <= 24'h0000ff;
		12'd0371: rd_data_1 <= 24'h0000ff;
		12'd0372: rd_data_1 <= 24'h0000ff;
		12'd0373: rd_data_1 <= 24'h0000ff;
		12'd0374: rd_data_1 <= 24'h0000ff;
		12'd0375: rd_data_1 <= 24'h0000ff;
		12'd0376: rd_data_1 <= 24'h000000;
		12'd0377: rd_data_1 <= 24'h000000;
		12'd0378: rd_data_1 <= 24'h000000;
		12'd0379: rd_data_1 <= 24'h000000;
		12'd0380: rd_data_1 <= 24'h000000;
		12'd0381: rd_data_1 <= 24'h000000;
		12'd0382: rd_data_1 <= 24'h000000;
		12'd0383: rd_data_1 <= 24'h000000;
		12'd0384: rd_data_1 <= 24'hffffff;
		12'd0385: rd_data_1 <= 24'hffffff;
		12'd0386: rd_data_1 <= 24'hffffff;
		12'd0387: rd_data_1 <= 24'hffffff;
		12'd0388: rd_data_1 <= 24'hffffff;
		12'd0389: rd_data_1 <= 24'hffffff;
		12'd0390: rd_data_1 <= 24'hffffff;
		12'd0391: rd_data_1 <= 24'hffffff;
		12'd0392: rd_data_1 <= 24'hffff00;
		12'd0393: rd_data_1 <= 24'hffff00;
		12'd0394: rd_data_1 <= 24'hffff00;
		12'd0395: rd_data_1 <= 24'hffff00;
		12'd0396: rd_data_1 <= 24'hffff00;
		12'd0397: rd_data_1 <= 24'hffff00;
		12'd0398: rd_data_1 <= 24'hffff00;
		12'd0399: rd_data_1 <= 24'hffff00;
		12'd0400: rd_data_1 <= 24'h00ffff;
		12'd0401: rd_data_1 <= 24'h00ffff;
		12'd0402: rd_data_1 <= 24'h00ffff;
		12'd0403: rd_data_1 <= 24'h00ffff;
		12'd0404: rd_data_1 <= 24'h00ffff;
		12'd0405: rd_data_1 <= 24'h00ffff;
		12'd0406: rd_data_1 <= 24'h00ffff;
		12'd0407: rd_data_1 <= 24'h00ffff;
		12'd0408: rd_data_1 <= 24'h00ff00;
		12'd0409: rd_data_1 <= 24'h00ff00;
		12'd0410: rd_data_1 <= 24'h00ff00;
		12'd0411: rd_data_1 <= 24'h00ff00;
		12'd0412: rd_data_1 <= 24'h00ff00;
		12'd0413: rd_data_1 <= 24'h00ff00;
		12'd0414: rd_data_1 <= 24'h00ff00;
		12'd0415: rd_data_1 <= 24'h00ff00;
		12'd0416: rd_data_1 <= 24'hff00ff;
		12'd0417: rd_data_1 <= 24'hff00ff;
		12'd0418: rd_data_1 <= 24'hff00ff;
		12'd0419: rd_data_1 <= 24'hff00ff;
		12'd0420: rd_data_1 <= 24'hff00ff;
		12'd0421: rd_data_1 <= 24'hff00ff;
		12'd0422: rd_data_1 <= 24'hff00ff;
		12'd0423: rd_data_1 <= 24'hff00ff;
		12'd0424: rd_data_1 <= 24'hff0000;
		12'd0425: rd_data_1 <= 24'hff0000;
		12'd0426: rd_data_1 <= 24'hff0000;
		12'd0427: rd_data_1 <= 24'hff0000;
		12'd0428: rd_data_1 <= 24'hff0000;
		12'd0429: rd_data_1 <= 24'hff0000;
		12'd0430: rd_data_1 <= 24'hff0000;
		12'd0431: rd_data_1 <= 24'hff0000;
		12'd0432: rd_data_1 <= 24'h0000ff;
		12'd0433: rd_data_1 <= 24'h0000ff;
		12'd0434: rd_data_1 <= 24'h0000ff;
		12'd0435: rd_data_1 <= 24'h0000ff;
		12'd0436: rd_data_1 <= 24'h0000ff;
		12'd0437: rd_data_1 <= 24'h0000ff;
		12'd0438: rd_data_1 <= 24'h0000ff;
		12'd0439: rd_data_1 <= 24'h0000ff;
		12'd0440: rd_data_1 <= 24'h000000;
		12'd0441: rd_data_1 <= 24'h000000;
		12'd0442: rd_data_1 <= 24'h000000;
		12'd0443: rd_data_1 <= 24'h000000;
		12'd0444: rd_data_1 <= 24'h000000;
		12'd0445: rd_data_1 <= 24'h000000;
		12'd0446: rd_data_1 <= 24'h000000;
		12'd0447: rd_data_1 <= 24'h000000;
		12'd0448: rd_data_1 <= 24'hffffff;
		12'd0449: rd_data_1 <= 24'hffffff;
		12'd0450: rd_data_1 <= 24'hffffff;
		12'd0451: rd_data_1 <= 24'hffffff;
		12'd0452: rd_data_1 <= 24'hffffff;
		12'd0453: rd_data_1 <= 24'hffffff;
		12'd0454: rd_data_1 <= 24'hffffff;
		12'd0455: rd_data_1 <= 24'hffffff;
		12'd0456: rd_data_1 <= 24'hffff00;
		12'd0457: rd_data_1 <= 24'hffff00;
		12'd0458: rd_data_1 <= 24'hffff00;
		12'd0459: rd_data_1 <= 24'hffff00;
		12'd0460: rd_data_1 <= 24'hffff00;
		12'd0461: rd_data_1 <= 24'hffff00;
		12'd0462: rd_data_1 <= 24'hffff00;
		12'd0463: rd_data_1 <= 24'hffff00;
		12'd0464: rd_data_1 <= 24'h00ffff;
		12'd0465: rd_data_1 <= 24'h00ffff;
		12'd0466: rd_data_1 <= 24'h00ffff;
		12'd0467: rd_data_1 <= 24'h00ffff;
		12'd0468: rd_data_1 <= 24'h00ffff;
		12'd0469: rd_data_1 <= 24'h00ffff;
		12'd0470: rd_data_1 <= 24'h00ffff;
		12'd0471: rd_data_1 <= 24'h00ffff;
		12'd0472: rd_data_1 <= 24'h00ff00;
		12'd0473: rd_data_1 <= 24'h00ff00;
		12'd0474: rd_data_1 <= 24'h00ff00;
		12'd0475: rd_data_1 <= 24'h00ff00;
		12'd0476: rd_data_1 <= 24'h00ff00;
		12'd0477: rd_data_1 <= 24'h00ff00;
		12'd0478: rd_data_1 <= 24'h00ff00;
		12'd0479: rd_data_1 <= 24'h00ff00;
		12'd0480: rd_data_1 <= 24'hff00ff;
		12'd0481: rd_data_1 <= 24'hff00ff;
		12'd0482: rd_data_1 <= 24'hff00ff;
		12'd0483: rd_data_1 <= 24'hff00ff;
		12'd0484: rd_data_1 <= 24'hff00ff;
		12'd0485: rd_data_1 <= 24'hff00ff;
		12'd0486: rd_data_1 <= 24'hff00ff;
		12'd0487: rd_data_1 <= 24'hff00ff;
		12'd0488: rd_data_1 <= 24'hff0000;
		12'd0489: rd_data_1 <= 24'hff0000;
		12'd0490: rd_data_1 <= 24'hff0000;
		12'd0491: rd_data_1 <= 24'hff0000;
		12'd0492: rd_data_1 <= 24'hff0000;
		12'd0493: rd_data_1 <= 24'hff0000;
		12'd0494: rd_data_1 <= 24'hff0000;
		12'd0495: rd_data_1 <= 24'hff0000;
		12'd0496: rd_data_1 <= 24'h0000ff;
		12'd0497: rd_data_1 <= 24'h0000ff;
		12'd0498: rd_data_1 <= 24'h0000ff;
		12'd0499: rd_data_1 <= 24'h0000ff;
		12'd0500: rd_data_1 <= 24'h0000ff;
		12'd0501: rd_data_1 <= 24'h0000ff;
		12'd0502: rd_data_1 <= 24'h0000ff;
		12'd0503: rd_data_1 <= 24'h0000ff;
		12'd0504: rd_data_1 <= 24'h000000;
		12'd0505: rd_data_1 <= 24'h000000;
		12'd0506: rd_data_1 <= 24'h000000;
		12'd0507: rd_data_1 <= 24'h000000;
		12'd0508: rd_data_1 <= 24'h000000;
		12'd0509: rd_data_1 <= 24'h000000;
		12'd0510: rd_data_1 <= 24'h000000;
		12'd0511: rd_data_1 <= 24'h000000;
		12'd0512: rd_data_1 <= 24'hffffff;
		12'd0513: rd_data_1 <= 24'hffffff;
		12'd0514: rd_data_1 <= 24'hffffff;
		12'd0515: rd_data_1 <= 24'hffffff;
		12'd0516: rd_data_1 <= 24'hffffff;
		12'd0517: rd_data_1 <= 24'hffffff;
		12'd0518: rd_data_1 <= 24'hffffff;
		12'd0519: rd_data_1 <= 24'hffffff;
		12'd0520: rd_data_1 <= 24'hffff00;
		12'd0521: rd_data_1 <= 24'hffff00;
		12'd0522: rd_data_1 <= 24'hffff00;
		12'd0523: rd_data_1 <= 24'hffff00;
		12'd0524: rd_data_1 <= 24'hffff00;
		12'd0525: rd_data_1 <= 24'hffff00;
		12'd0526: rd_data_1 <= 24'hffff00;
		12'd0527: rd_data_1 <= 24'hffff00;
		12'd0528: rd_data_1 <= 24'h00ffff;
		12'd0529: rd_data_1 <= 24'h00ffff;
		12'd0530: rd_data_1 <= 24'h00ffff;
		12'd0531: rd_data_1 <= 24'h00ffff;
		12'd0532: rd_data_1 <= 24'h00ffff;
		12'd0533: rd_data_1 <= 24'h00ffff;
		12'd0534: rd_data_1 <= 24'h00ffff;
		12'd0535: rd_data_1 <= 24'h00ffff;
		12'd0536: rd_data_1 <= 24'h00ff00;
		12'd0537: rd_data_1 <= 24'h00ff00;
		12'd0538: rd_data_1 <= 24'h00ff00;
		12'd0539: rd_data_1 <= 24'h00ff00;
		12'd0540: rd_data_1 <= 24'h00ff00;
		12'd0541: rd_data_1 <= 24'h00ff00;
		12'd0542: rd_data_1 <= 24'h00ff00;
		12'd0543: rd_data_1 <= 24'h00ff00;
		12'd0544: rd_data_1 <= 24'hff00ff;
		12'd0545: rd_data_1 <= 24'hff00ff;
		12'd0546: rd_data_1 <= 24'hff00ff;
		12'd0547: rd_data_1 <= 24'hff00ff;
		12'd0548: rd_data_1 <= 24'hff00ff;
		12'd0549: rd_data_1 <= 24'hff00ff;
		12'd0550: rd_data_1 <= 24'hff00ff;
		12'd0551: rd_data_1 <= 24'hff00ff;
		12'd0552: rd_data_1 <= 24'hff0000;
		12'd0553: rd_data_1 <= 24'hff0000;
		12'd0554: rd_data_1 <= 24'hff0000;
		12'd0555: rd_data_1 <= 24'hff0000;
		12'd0556: rd_data_1 <= 24'hff0000;
		12'd0557: rd_data_1 <= 24'hff0000;
		12'd0558: rd_data_1 <= 24'hff0000;
		12'd0559: rd_data_1 <= 24'hff0000;
		12'd0560: rd_data_1 <= 24'h0000ff;
		12'd0561: rd_data_1 <= 24'h0000ff;
		12'd0562: rd_data_1 <= 24'h0000ff;
		12'd0563: rd_data_1 <= 24'h0000ff;
		12'd0564: rd_data_1 <= 24'h0000ff;
		12'd0565: rd_data_1 <= 24'h0000ff;
		12'd0566: rd_data_1 <= 24'h0000ff;
		12'd0567: rd_data_1 <= 24'h0000ff;
		12'd0568: rd_data_1 <= 24'h000000;
		12'd0569: rd_data_1 <= 24'h000000;
		12'd0570: rd_data_1 <= 24'h000000;
		12'd0571: rd_data_1 <= 24'h000000;
		12'd0572: rd_data_1 <= 24'h000000;
		12'd0573: rd_data_1 <= 24'h000000;
		12'd0574: rd_data_1 <= 24'h000000;
		12'd0575: rd_data_1 <= 24'h000000;
		12'd0576: rd_data_1 <= 24'hffffff;
		12'd0577: rd_data_1 <= 24'hffffff;
		12'd0578: rd_data_1 <= 24'hffffff;
		12'd0579: rd_data_1 <= 24'hffffff;
		12'd0580: rd_data_1 <= 24'hffffff;
		12'd0581: rd_data_1 <= 24'hffffff;
		12'd0582: rd_data_1 <= 24'hffffff;
		12'd0583: rd_data_1 <= 24'hffffff;
		12'd0584: rd_data_1 <= 24'hffff00;
		12'd0585: rd_data_1 <= 24'hffff00;
		12'd0586: rd_data_1 <= 24'hffff00;
		12'd0587: rd_data_1 <= 24'hffff00;
		12'd0588: rd_data_1 <= 24'hffff00;
		12'd0589: rd_data_1 <= 24'hffff00;
		12'd0590: rd_data_1 <= 24'hffff00;
		12'd0591: rd_data_1 <= 24'hffff00;
		12'd0592: rd_data_1 <= 24'h00ffff;
		12'd0593: rd_data_1 <= 24'h00ffff;
		12'd0594: rd_data_1 <= 24'h00ffff;
		12'd0595: rd_data_1 <= 24'h00ffff;
		12'd0596: rd_data_1 <= 24'h00ffff;
		12'd0597: rd_data_1 <= 24'h00ffff;
		12'd0598: rd_data_1 <= 24'h00ffff;
		12'd0599: rd_data_1 <= 24'h00ffff;
		12'd0600: rd_data_1 <= 24'h00ff00;
		12'd0601: rd_data_1 <= 24'h00ff00;
		12'd0602: rd_data_1 <= 24'h00ff00;
		12'd0603: rd_data_1 <= 24'h00ff00;
		12'd0604: rd_data_1 <= 24'h00ff00;
		12'd0605: rd_data_1 <= 24'h00ff00;
		12'd0606: rd_data_1 <= 24'h00ff00;
		12'd0607: rd_data_1 <= 24'h00ff00;
		12'd0608: rd_data_1 <= 24'hff00ff;
		12'd0609: rd_data_1 <= 24'hff00ff;
		12'd0610: rd_data_1 <= 24'hff00ff;
		12'd0611: rd_data_1 <= 24'hff00ff;
		12'd0612: rd_data_1 <= 24'hff00ff;
		12'd0613: rd_data_1 <= 24'hff00ff;
		12'd0614: rd_data_1 <= 24'hff00ff;
		12'd0615: rd_data_1 <= 24'hff00ff;
		12'd0616: rd_data_1 <= 24'hff0000;
		12'd0617: rd_data_1 <= 24'hff0000;
		12'd0618: rd_data_1 <= 24'hff0000;
		12'd0619: rd_data_1 <= 24'hff0000;
		12'd0620: rd_data_1 <= 24'hff0000;
		12'd0621: rd_data_1 <= 24'hff0000;
		12'd0622: rd_data_1 <= 24'hff0000;
		12'd0623: rd_data_1 <= 24'hff0000;
		12'd0624: rd_data_1 <= 24'h0000ff;
		12'd0625: rd_data_1 <= 24'h0000ff;
		12'd0626: rd_data_1 <= 24'h0000ff;
		12'd0627: rd_data_1 <= 24'h0000ff;
		12'd0628: rd_data_1 <= 24'h0000ff;
		12'd0629: rd_data_1 <= 24'h0000ff;
		12'd0630: rd_data_1 <= 24'h0000ff;
		12'd0631: rd_data_1 <= 24'h0000ff;
		12'd0632: rd_data_1 <= 24'h000000;
		12'd0633: rd_data_1 <= 24'h000000;
		12'd0634: rd_data_1 <= 24'h000000;
		12'd0635: rd_data_1 <= 24'h000000;
		12'd0636: rd_data_1 <= 24'h000000;
		12'd0637: rd_data_1 <= 24'h000000;
		12'd0638: rd_data_1 <= 24'h000000;
		12'd0639: rd_data_1 <= 24'h000000;
		12'd0640: rd_data_1 <= 24'hffffff;
		12'd0641: rd_data_1 <= 24'hffffff;
		12'd0642: rd_data_1 <= 24'hffffff;
		12'd0643: rd_data_1 <= 24'hffffff;
		12'd0644: rd_data_1 <= 24'hffffff;
		12'd0645: rd_data_1 <= 24'hffffff;
		12'd0646: rd_data_1 <= 24'hffffff;
		12'd0647: rd_data_1 <= 24'hffffff;
		12'd0648: rd_data_1 <= 24'hffff00;
		12'd0649: rd_data_1 <= 24'hffff00;
		12'd0650: rd_data_1 <= 24'hffff00;
		12'd0651: rd_data_1 <= 24'hffff00;
		12'd0652: rd_data_1 <= 24'hffff00;
		12'd0653: rd_data_1 <= 24'hffff00;
		12'd0654: rd_data_1 <= 24'hffff00;
		12'd0655: rd_data_1 <= 24'hffff00;
		12'd0656: rd_data_1 <= 24'h00ffff;
		12'd0657: rd_data_1 <= 24'h00ffff;
		12'd0658: rd_data_1 <= 24'h00ffff;
		12'd0659: rd_data_1 <= 24'h00ffff;
		12'd0660: rd_data_1 <= 24'h00ffff;
		12'd0661: rd_data_1 <= 24'h00ffff;
		12'd0662: rd_data_1 <= 24'h00ffff;
		12'd0663: rd_data_1 <= 24'h00ffff;
		12'd0664: rd_data_1 <= 24'h00ff00;
		12'd0665: rd_data_1 <= 24'h00ff00;
		12'd0666: rd_data_1 <= 24'h00ff00;
		12'd0667: rd_data_1 <= 24'h00ff00;
		12'd0668: rd_data_1 <= 24'h00ff00;
		12'd0669: rd_data_1 <= 24'h00ff00;
		12'd0670: rd_data_1 <= 24'h00ff00;
		12'd0671: rd_data_1 <= 24'h00ff00;
		12'd0672: rd_data_1 <= 24'hff00ff;
		12'd0673: rd_data_1 <= 24'hff00ff;
		12'd0674: rd_data_1 <= 24'hff00ff;
		12'd0675: rd_data_1 <= 24'hff00ff;
		12'd0676: rd_data_1 <= 24'hff00ff;
		12'd0677: rd_data_1 <= 24'hff00ff;
		12'd0678: rd_data_1 <= 24'hff00ff;
		12'd0679: rd_data_1 <= 24'hff00ff;
		12'd0680: rd_data_1 <= 24'hff0000;
		12'd0681: rd_data_1 <= 24'hff0000;
		12'd0682: rd_data_1 <= 24'hff0000;
		12'd0683: rd_data_1 <= 24'hff0000;
		12'd0684: rd_data_1 <= 24'hff0000;
		12'd0685: rd_data_1 <= 24'hff0000;
		12'd0686: rd_data_1 <= 24'hff0000;
		12'd0687: rd_data_1 <= 24'hff0000;
		12'd0688: rd_data_1 <= 24'h0000ff;
		12'd0689: rd_data_1 <= 24'h0000ff;
		12'd0690: rd_data_1 <= 24'h0000ff;
		12'd0691: rd_data_1 <= 24'h0000ff;
		12'd0692: rd_data_1 <= 24'h0000ff;
		12'd0693: rd_data_1 <= 24'h0000ff;
		12'd0694: rd_data_1 <= 24'h0000ff;
		12'd0695: rd_data_1 <= 24'h0000ff;
		12'd0696: rd_data_1 <= 24'h000000;
		12'd0697: rd_data_1 <= 24'h000000;
		12'd0698: rd_data_1 <= 24'h000000;
		12'd0699: rd_data_1 <= 24'h000000;
		12'd0700: rd_data_1 <= 24'h000000;
		12'd0701: rd_data_1 <= 24'h000000;
		12'd0702: rd_data_1 <= 24'h000000;
		12'd0703: rd_data_1 <= 24'h000000;
		12'd0704: rd_data_1 <= 24'hffffff;
		12'd0705: rd_data_1 <= 24'hffffff;
		12'd0706: rd_data_1 <= 24'hffffff;
		12'd0707: rd_data_1 <= 24'hffffff;
		12'd0708: rd_data_1 <= 24'hffffff;
		12'd0709: rd_data_1 <= 24'hffffff;
		12'd0710: rd_data_1 <= 24'hffffff;
		12'd0711: rd_data_1 <= 24'hffffff;
		12'd0712: rd_data_1 <= 24'hffff00;
		12'd0713: rd_data_1 <= 24'hffff00;
		12'd0714: rd_data_1 <= 24'hffff00;
		12'd0715: rd_data_1 <= 24'hffff00;
		12'd0716: rd_data_1 <= 24'hffff00;
		12'd0717: rd_data_1 <= 24'hffff00;
		12'd0718: rd_data_1 <= 24'hffff00;
		12'd0719: rd_data_1 <= 24'hffff00;
		12'd0720: rd_data_1 <= 24'h00ffff;
		12'd0721: rd_data_1 <= 24'h00ffff;
		12'd0722: rd_data_1 <= 24'h00ffff;
		12'd0723: rd_data_1 <= 24'h00ffff;
		12'd0724: rd_data_1 <= 24'h00ffff;
		12'd0725: rd_data_1 <= 24'h00ffff;
		12'd0726: rd_data_1 <= 24'h00ffff;
		12'd0727: rd_data_1 <= 24'h00ffff;
		12'd0728: rd_data_1 <= 24'h00ff00;
		12'd0729: rd_data_1 <= 24'h00ff00;
		12'd0730: rd_data_1 <= 24'h00ff00;
		12'd0731: rd_data_1 <= 24'h00ff00;
		12'd0732: rd_data_1 <= 24'h00ff00;
		12'd0733: rd_data_1 <= 24'h00ff00;
		12'd0734: rd_data_1 <= 24'h00ff00;
		12'd0735: rd_data_1 <= 24'h00ff00;
		12'd0736: rd_data_1 <= 24'hff00ff;
		12'd0737: rd_data_1 <= 24'hff00ff;
		12'd0738: rd_data_1 <= 24'hff00ff;
		12'd0739: rd_data_1 <= 24'hff00ff;
		12'd0740: rd_data_1 <= 24'hff00ff;
		12'd0741: rd_data_1 <= 24'hff00ff;
		12'd0742: rd_data_1 <= 24'hff00ff;
		12'd0743: rd_data_1 <= 24'hff00ff;
		12'd0744: rd_data_1 <= 24'hff0000;
		12'd0745: rd_data_1 <= 24'hff0000;
		12'd0746: rd_data_1 <= 24'hff0000;
		12'd0747: rd_data_1 <= 24'hff0000;
		12'd0748: rd_data_1 <= 24'hff0000;
		12'd0749: rd_data_1 <= 24'hff0000;
		12'd0750: rd_data_1 <= 24'hff0000;
		12'd0751: rd_data_1 <= 24'hff0000;
		12'd0752: rd_data_1 <= 24'h0000ff;
		12'd0753: rd_data_1 <= 24'h0000ff;
		12'd0754: rd_data_1 <= 24'h0000ff;
		12'd0755: rd_data_1 <= 24'h0000ff;
		12'd0756: rd_data_1 <= 24'h0000ff;
		12'd0757: rd_data_1 <= 24'h0000ff;
		12'd0758: rd_data_1 <= 24'h0000ff;
		12'd0759: rd_data_1 <= 24'h0000ff;
		12'd0760: rd_data_1 <= 24'h000000;
		12'd0761: rd_data_1 <= 24'h000000;
		12'd0762: rd_data_1 <= 24'h000000;
		12'd0763: rd_data_1 <= 24'h000000;
		12'd0764: rd_data_1 <= 24'h000000;
		12'd0765: rd_data_1 <= 24'h000000;
		12'd0766: rd_data_1 <= 24'h000000;
		12'd0767: rd_data_1 <= 24'h000000;
		12'd0768: rd_data_1 <= 24'hffffff;
		12'd0769: rd_data_1 <= 24'hffffff;
		12'd0770: rd_data_1 <= 24'hffffff;
		12'd0771: rd_data_1 <= 24'hffffff;
		12'd0772: rd_data_1 <= 24'hffffff;
		12'd0773: rd_data_1 <= 24'hffffff;
		12'd0774: rd_data_1 <= 24'hffffff;
		12'd0775: rd_data_1 <= 24'hffffff;
		12'd0776: rd_data_1 <= 24'hffff00;
		12'd0777: rd_data_1 <= 24'hffff00;
		12'd0778: rd_data_1 <= 24'hffff00;
		12'd0779: rd_data_1 <= 24'hffff00;
		12'd0780: rd_data_1 <= 24'hffff00;
		12'd0781: rd_data_1 <= 24'hffff00;
		12'd0782: rd_data_1 <= 24'hffff00;
		12'd0783: rd_data_1 <= 24'hffff00;
		12'd0784: rd_data_1 <= 24'h00ffff;
		12'd0785: rd_data_1 <= 24'h00ffff;
		12'd0786: rd_data_1 <= 24'h00ffff;
		12'd0787: rd_data_1 <= 24'h00ffff;
		12'd0788: rd_data_1 <= 24'h00ffff;
		12'd0789: rd_data_1 <= 24'h00ffff;
		12'd0790: rd_data_1 <= 24'h00ffff;
		12'd0791: rd_data_1 <= 24'h00ffff;
		12'd0792: rd_data_1 <= 24'h00ff00;
		12'd0793: rd_data_1 <= 24'h00ff00;
		12'd0794: rd_data_1 <= 24'h00ff00;
		12'd0795: rd_data_1 <= 24'h00ff00;
		12'd0796: rd_data_1 <= 24'h00ff00;
		12'd0797: rd_data_1 <= 24'h00ff00;
		12'd0798: rd_data_1 <= 24'h00ff00;
		12'd0799: rd_data_1 <= 24'h00ff00;
		12'd0800: rd_data_1 <= 24'hff00ff;
		12'd0801: rd_data_1 <= 24'hff00ff;
		12'd0802: rd_data_1 <= 24'hff00ff;
		12'd0803: rd_data_1 <= 24'hff00ff;
		12'd0804: rd_data_1 <= 24'hff00ff;
		12'd0805: rd_data_1 <= 24'hff00ff;
		12'd0806: rd_data_1 <= 24'hff00ff;
		12'd0807: rd_data_1 <= 24'hff00ff;
		12'd0808: rd_data_1 <= 24'hff0000;
		12'd0809: rd_data_1 <= 24'hff0000;
		12'd0810: rd_data_1 <= 24'hff0000;
		12'd0811: rd_data_1 <= 24'hff0000;
		12'd0812: rd_data_1 <= 24'hff0000;
		12'd0813: rd_data_1 <= 24'hff0000;
		12'd0814: rd_data_1 <= 24'hff0000;
		12'd0815: rd_data_1 <= 24'hff0000;
		12'd0816: rd_data_1 <= 24'h0000ff;
		12'd0817: rd_data_1 <= 24'h0000ff;
		12'd0818: rd_data_1 <= 24'h0000ff;
		12'd0819: rd_data_1 <= 24'h0000ff;
		12'd0820: rd_data_1 <= 24'h0000ff;
		12'd0821: rd_data_1 <= 24'h0000ff;
		12'd0822: rd_data_1 <= 24'h0000ff;
		12'd0823: rd_data_1 <= 24'h0000ff;
		12'd0824: rd_data_1 <= 24'h000000;
		12'd0825: rd_data_1 <= 24'h000000;
		12'd0826: rd_data_1 <= 24'h000000;
		12'd0827: rd_data_1 <= 24'h000000;
		12'd0828: rd_data_1 <= 24'h000000;
		12'd0829: rd_data_1 <= 24'h000000;
		12'd0830: rd_data_1 <= 24'h000000;
		12'd0831: rd_data_1 <= 24'h000000;
		12'd0832: rd_data_1 <= 24'hffffff;
		12'd0833: rd_data_1 <= 24'hffffff;
		12'd0834: rd_data_1 <= 24'hffffff;
		12'd0835: rd_data_1 <= 24'hffffff;
		12'd0836: rd_data_1 <= 24'hffffff;
		12'd0837: rd_data_1 <= 24'hffffff;
		12'd0838: rd_data_1 <= 24'hffffff;
		12'd0839: rd_data_1 <= 24'hffffff;
		12'd0840: rd_data_1 <= 24'hffff00;
		12'd0841: rd_data_1 <= 24'hffff00;
		12'd0842: rd_data_1 <= 24'hffff00;
		12'd0843: rd_data_1 <= 24'hffff00;
		12'd0844: rd_data_1 <= 24'hffff00;
		12'd0845: rd_data_1 <= 24'hffff00;
		12'd0846: rd_data_1 <= 24'hffff00;
		12'd0847: rd_data_1 <= 24'hffff00;
		12'd0848: rd_data_1 <= 24'h00ffff;
		12'd0849: rd_data_1 <= 24'h00ffff;
		12'd0850: rd_data_1 <= 24'h00ffff;
		12'd0851: rd_data_1 <= 24'h00ffff;
		12'd0852: rd_data_1 <= 24'h00ffff;
		12'd0853: rd_data_1 <= 24'h00ffff;
		12'd0854: rd_data_1 <= 24'h00ffff;
		12'd0855: rd_data_1 <= 24'h00ffff;
		12'd0856: rd_data_1 <= 24'h00ff00;
		12'd0857: rd_data_1 <= 24'h00ff00;
		12'd0858: rd_data_1 <= 24'h00ff00;
		12'd0859: rd_data_1 <= 24'h00ff00;
		12'd0860: rd_data_1 <= 24'h00ff00;
		12'd0861: rd_data_1 <= 24'h00ff00;
		12'd0862: rd_data_1 <= 24'h00ff00;
		12'd0863: rd_data_1 <= 24'h00ff00;
		12'd0864: rd_data_1 <= 24'hff00ff;
		12'd0865: rd_data_1 <= 24'hff00ff;
		12'd0866: rd_data_1 <= 24'hff00ff;
		12'd0867: rd_data_1 <= 24'hff00ff;
		12'd0868: rd_data_1 <= 24'hff00ff;
		12'd0869: rd_data_1 <= 24'hff00ff;
		12'd0870: rd_data_1 <= 24'hff00ff;
		12'd0871: rd_data_1 <= 24'hff00ff;
		12'd0872: rd_data_1 <= 24'hff0000;
		12'd0873: rd_data_1 <= 24'hff0000;
		12'd0874: rd_data_1 <= 24'hff0000;
		12'd0875: rd_data_1 <= 24'hff0000;
		12'd0876: rd_data_1 <= 24'hff0000;
		12'd0877: rd_data_1 <= 24'hff0000;
		12'd0878: rd_data_1 <= 24'hff0000;
		12'd0879: rd_data_1 <= 24'hff0000;
		12'd0880: rd_data_1 <= 24'h0000ff;
		12'd0881: rd_data_1 <= 24'h0000ff;
		12'd0882: rd_data_1 <= 24'h0000ff;
		12'd0883: rd_data_1 <= 24'h0000ff;
		12'd0884: rd_data_1 <= 24'h0000ff;
		12'd0885: rd_data_1 <= 24'h0000ff;
		12'd0886: rd_data_1 <= 24'h0000ff;
		12'd0887: rd_data_1 <= 24'h0000ff;
		12'd0888: rd_data_1 <= 24'h000000;
		12'd0889: rd_data_1 <= 24'h000000;
		12'd0890: rd_data_1 <= 24'h000000;
		12'd0891: rd_data_1 <= 24'h000000;
		12'd0892: rd_data_1 <= 24'h000000;
		12'd0893: rd_data_1 <= 24'h000000;
		12'd0894: rd_data_1 <= 24'h000000;
		12'd0895: rd_data_1 <= 24'h000000;
		12'd0896: rd_data_1 <= 24'hffffff;
		12'd0897: rd_data_1 <= 24'hffffff;
		12'd0898: rd_data_1 <= 24'hffffff;
		12'd0899: rd_data_1 <= 24'hffffff;
		12'd0900: rd_data_1 <= 24'hffffff;
		12'd0901: rd_data_1 <= 24'hffffff;
		12'd0902: rd_data_1 <= 24'hffffff;
		12'd0903: rd_data_1 <= 24'hffffff;
		12'd0904: rd_data_1 <= 24'hffff00;
		12'd0905: rd_data_1 <= 24'hffff00;
		12'd0906: rd_data_1 <= 24'hffff00;
		12'd0907: rd_data_1 <= 24'hffff00;
		12'd0908: rd_data_1 <= 24'hffff00;
		12'd0909: rd_data_1 <= 24'hffff00;
		12'd0910: rd_data_1 <= 24'hffff00;
		12'd0911: rd_data_1 <= 24'hffff00;
		12'd0912: rd_data_1 <= 24'h00ffff;
		12'd0913: rd_data_1 <= 24'h00ffff;
		12'd0914: rd_data_1 <= 24'h00ffff;
		12'd0915: rd_data_1 <= 24'h00ffff;
		12'd0916: rd_data_1 <= 24'h00ffff;
		12'd0917: rd_data_1 <= 24'h00ffff;
		12'd0918: rd_data_1 <= 24'h00ffff;
		12'd0919: rd_data_1 <= 24'h00ffff;
		12'd0920: rd_data_1 <= 24'h00ff00;
		12'd0921: rd_data_1 <= 24'h00ff00;
		12'd0922: rd_data_1 <= 24'h00ff00;
		12'd0923: rd_data_1 <= 24'h00ff00;
		12'd0924: rd_data_1 <= 24'h00ff00;
		12'd0925: rd_data_1 <= 24'h00ff00;
		12'd0926: rd_data_1 <= 24'h00ff00;
		12'd0927: rd_data_1 <= 24'h00ff00;
		12'd0928: rd_data_1 <= 24'hff00ff;
		12'd0929: rd_data_1 <= 24'hff00ff;
		12'd0930: rd_data_1 <= 24'hff00ff;
		12'd0931: rd_data_1 <= 24'hff00ff;
		12'd0932: rd_data_1 <= 24'hff00ff;
		12'd0933: rd_data_1 <= 24'hff00ff;
		12'd0934: rd_data_1 <= 24'hff00ff;
		12'd0935: rd_data_1 <= 24'hff00ff;
		12'd0936: rd_data_1 <= 24'hff0000;
		12'd0937: rd_data_1 <= 24'hff0000;
		12'd0938: rd_data_1 <= 24'hff0000;
		12'd0939: rd_data_1 <= 24'hff0000;
		12'd0940: rd_data_1 <= 24'hff0000;
		12'd0941: rd_data_1 <= 24'hff0000;
		12'd0942: rd_data_1 <= 24'hff0000;
		12'd0943: rd_data_1 <= 24'hff0000;
		12'd0944: rd_data_1 <= 24'h0000ff;
		12'd0945: rd_data_1 <= 24'h0000ff;
		12'd0946: rd_data_1 <= 24'h0000ff;
		12'd0947: rd_data_1 <= 24'h0000ff;
		12'd0948: rd_data_1 <= 24'h0000ff;
		12'd0949: rd_data_1 <= 24'h0000ff;
		12'd0950: rd_data_1 <= 24'h0000ff;
		12'd0951: rd_data_1 <= 24'h0000ff;
		12'd0952: rd_data_1 <= 24'h000000;
		12'd0953: rd_data_1 <= 24'h000000;
		12'd0954: rd_data_1 <= 24'h000000;
		12'd0955: rd_data_1 <= 24'h000000;
		12'd0956: rd_data_1 <= 24'h000000;
		12'd0957: rd_data_1 <= 24'h000000;
		12'd0958: rd_data_1 <= 24'h000000;
		12'd0959: rd_data_1 <= 24'h000000;
		12'd0960: rd_data_1 <= 24'hffffff;
		12'd0961: rd_data_1 <= 24'hffffff;
		12'd0962: rd_data_1 <= 24'hffffff;
		12'd0963: rd_data_1 <= 24'hffffff;
		12'd0964: rd_data_1 <= 24'hffffff;
		12'd0965: rd_data_1 <= 24'hffffff;
		12'd0966: rd_data_1 <= 24'hffffff;
		12'd0967: rd_data_1 <= 24'hffffff;
		12'd0968: rd_data_1 <= 24'hffff00;
		12'd0969: rd_data_1 <= 24'hffff00;
		12'd0970: rd_data_1 <= 24'hffff00;
		12'd0971: rd_data_1 <= 24'hffff00;
		12'd0972: rd_data_1 <= 24'hffff00;
		12'd0973: rd_data_1 <= 24'hffff00;
		12'd0974: rd_data_1 <= 24'hffff00;
		12'd0975: rd_data_1 <= 24'hffff00;
		12'd0976: rd_data_1 <= 24'h00ffff;
		12'd0977: rd_data_1 <= 24'h00ffff;
		12'd0978: rd_data_1 <= 24'h00ffff;
		12'd0979: rd_data_1 <= 24'h00ffff;
		12'd0980: rd_data_1 <= 24'h00ffff;
		12'd0981: rd_data_1 <= 24'h00ffff;
		12'd0982: rd_data_1 <= 24'h00ffff;
		12'd0983: rd_data_1 <= 24'h00ffff;
		12'd0984: rd_data_1 <= 24'h00ff00;
		12'd0985: rd_data_1 <= 24'h00ff00;
		12'd0986: rd_data_1 <= 24'h00ff00;
		12'd0987: rd_data_1 <= 24'h00ff00;
		12'd0988: rd_data_1 <= 24'h00ff00;
		12'd0989: rd_data_1 <= 24'h00ff00;
		12'd0990: rd_data_1 <= 24'h00ff00;
		12'd0991: rd_data_1 <= 24'h00ff00;
		12'd0992: rd_data_1 <= 24'hff00ff;
		12'd0993: rd_data_1 <= 24'hff00ff;
		12'd0994: rd_data_1 <= 24'hff00ff;
		12'd0995: rd_data_1 <= 24'hff00ff;
		12'd0996: rd_data_1 <= 24'hff00ff;
		12'd0997: rd_data_1 <= 24'hff00ff;
		12'd0998: rd_data_1 <= 24'hff00ff;
		12'd0999: rd_data_1 <= 24'hff00ff;
		12'd1000: rd_data_1 <= 24'hff0000;
		12'd1001: rd_data_1 <= 24'hff0000;
		12'd1002: rd_data_1 <= 24'hff0000;
		12'd1003: rd_data_1 <= 24'hff0000;
		12'd1004: rd_data_1 <= 24'hff0000;
		12'd1005: rd_data_1 <= 24'hff0000;
		12'd1006: rd_data_1 <= 24'hff0000;
		12'd1007: rd_data_1 <= 24'hff0000;
		12'd1008: rd_data_1 <= 24'h0000ff;
		12'd1009: rd_data_1 <= 24'h0000ff;
		12'd1010: rd_data_1 <= 24'h0000ff;
		12'd1011: rd_data_1 <= 24'h0000ff;
		12'd1012: rd_data_1 <= 24'h0000ff;
		12'd1013: rd_data_1 <= 24'h0000ff;
		12'd1014: rd_data_1 <= 24'h0000ff;
		12'd1015: rd_data_1 <= 24'h0000ff;
		12'd1016: rd_data_1 <= 24'h000000;
		12'd1017: rd_data_1 <= 24'h000000;
		12'd1018: rd_data_1 <= 24'h000000;
		12'd1019: rd_data_1 <= 24'h000000;
		12'd1020: rd_data_1 <= 24'h000000;
		12'd1021: rd_data_1 <= 24'h000000;
		12'd1022: rd_data_1 <= 24'h000000;
		12'd1023: rd_data_1 <= 24'h000000;
		12'd1024: rd_data_1 <= 24'hffffff;
		12'd1025: rd_data_1 <= 24'hffffff;
		12'd1026: rd_data_1 <= 24'hffffff;
		12'd1027: rd_data_1 <= 24'hffffff;
		12'd1028: rd_data_1 <= 24'hffffff;
		12'd1029: rd_data_1 <= 24'hffffff;
		12'd1030: rd_data_1 <= 24'hffffff;
		12'd1031: rd_data_1 <= 24'hffffff;
		12'd1032: rd_data_1 <= 24'hffff00;
		12'd1033: rd_data_1 <= 24'hffff00;
		12'd1034: rd_data_1 <= 24'hffff00;
		12'd1035: rd_data_1 <= 24'hffff00;
		12'd1036: rd_data_1 <= 24'hffff00;
		12'd1037: rd_data_1 <= 24'hffff00;
		12'd1038: rd_data_1 <= 24'hffff00;
		12'd1039: rd_data_1 <= 24'hffff00;
		12'd1040: rd_data_1 <= 24'h00ffff;
		12'd1041: rd_data_1 <= 24'h00ffff;
		12'd1042: rd_data_1 <= 24'h00ffff;
		12'd1043: rd_data_1 <= 24'h00ffff;
		12'd1044: rd_data_1 <= 24'h00ffff;
		12'd1045: rd_data_1 <= 24'h00ffff;
		12'd1046: rd_data_1 <= 24'h00ffff;
		12'd1047: rd_data_1 <= 24'h00ffff;
		12'd1048: rd_data_1 <= 24'h00ff00;
		12'd1049: rd_data_1 <= 24'h00ff00;
		12'd1050: rd_data_1 <= 24'h00ff00;
		12'd1051: rd_data_1 <= 24'h00ff00;
		12'd1052: rd_data_1 <= 24'h00ff00;
		12'd1053: rd_data_1 <= 24'h00ff00;
		12'd1054: rd_data_1 <= 24'h00ff00;
		12'd1055: rd_data_1 <= 24'h00ff00;
		12'd1056: rd_data_1 <= 24'hff00ff;
		12'd1057: rd_data_1 <= 24'hff00ff;
		12'd1058: rd_data_1 <= 24'hff00ff;
		12'd1059: rd_data_1 <= 24'hff00ff;
		12'd1060: rd_data_1 <= 24'hff00ff;
		12'd1061: rd_data_1 <= 24'hff00ff;
		12'd1062: rd_data_1 <= 24'hff00ff;
		12'd1063: rd_data_1 <= 24'hff00ff;
		12'd1064: rd_data_1 <= 24'hff0000;
		12'd1065: rd_data_1 <= 24'hff0000;
		12'd1066: rd_data_1 <= 24'hff0000;
		12'd1067: rd_data_1 <= 24'hff0000;
		12'd1068: rd_data_1 <= 24'hff0000;
		12'd1069: rd_data_1 <= 24'hff0000;
		12'd1070: rd_data_1 <= 24'hff0000;
		12'd1071: rd_data_1 <= 24'hff0000;
		12'd1072: rd_data_1 <= 24'h0000ff;
		12'd1073: rd_data_1 <= 24'h0000ff;
		12'd1074: rd_data_1 <= 24'h0000ff;
		12'd1075: rd_data_1 <= 24'h0000ff;
		12'd1076: rd_data_1 <= 24'h0000ff;
		12'd1077: rd_data_1 <= 24'h0000ff;
		12'd1078: rd_data_1 <= 24'h0000ff;
		12'd1079: rd_data_1 <= 24'h0000ff;
		12'd1080: rd_data_1 <= 24'h000000;
		12'd1081: rd_data_1 <= 24'h000000;
		12'd1082: rd_data_1 <= 24'h000000;
		12'd1083: rd_data_1 <= 24'h000000;
		12'd1084: rd_data_1 <= 24'h000000;
		12'd1085: rd_data_1 <= 24'h000000;
		12'd1086: rd_data_1 <= 24'h000000;
		12'd1087: rd_data_1 <= 24'h000000;
		12'd1088: rd_data_1 <= 24'hffffff;
		12'd1089: rd_data_1 <= 24'hffffff;
		12'd1090: rd_data_1 <= 24'hffffff;
		12'd1091: rd_data_1 <= 24'hffffff;
		12'd1092: rd_data_1 <= 24'hffffff;
		12'd1093: rd_data_1 <= 24'hffffff;
		12'd1094: rd_data_1 <= 24'hffffff;
		12'd1095: rd_data_1 <= 24'hffffff;
		12'd1096: rd_data_1 <= 24'hffff00;
		12'd1097: rd_data_1 <= 24'hffff00;
		12'd1098: rd_data_1 <= 24'hffff00;
		12'd1099: rd_data_1 <= 24'hffff00;
		12'd1100: rd_data_1 <= 24'hffff00;
		12'd1101: rd_data_1 <= 24'hffff00;
		12'd1102: rd_data_1 <= 24'hffff00;
		12'd1103: rd_data_1 <= 24'hffff00;
		12'd1104: rd_data_1 <= 24'h00ffff;
		12'd1105: rd_data_1 <= 24'h00ffff;
		12'd1106: rd_data_1 <= 24'h00ffff;
		12'd1107: rd_data_1 <= 24'h00ffff;
		12'd1108: rd_data_1 <= 24'h00ffff;
		12'd1109: rd_data_1 <= 24'h00ffff;
		12'd1110: rd_data_1 <= 24'h00ffff;
		12'd1111: rd_data_1 <= 24'h00ffff;
		12'd1112: rd_data_1 <= 24'h00ff00;
		12'd1113: rd_data_1 <= 24'h00ff00;
		12'd1114: rd_data_1 <= 24'h00ff00;
		12'd1115: rd_data_1 <= 24'h00ff00;
		12'd1116: rd_data_1 <= 24'h00ff00;
		12'd1117: rd_data_1 <= 24'h00ff00;
		12'd1118: rd_data_1 <= 24'h00ff00;
		12'd1119: rd_data_1 <= 24'h00ff00;
		12'd1120: rd_data_1 <= 24'hff00ff;
		12'd1121: rd_data_1 <= 24'hff00ff;
		12'd1122: rd_data_1 <= 24'hff00ff;
		12'd1123: rd_data_1 <= 24'hff00ff;
		12'd1124: rd_data_1 <= 24'hff00ff;
		12'd1125: rd_data_1 <= 24'hff00ff;
		12'd1126: rd_data_1 <= 24'hff00ff;
		12'd1127: rd_data_1 <= 24'hff00ff;
		12'd1128: rd_data_1 <= 24'hff0000;
		12'd1129: rd_data_1 <= 24'hff0000;
		12'd1130: rd_data_1 <= 24'hff0000;
		12'd1131: rd_data_1 <= 24'hff0000;
		12'd1132: rd_data_1 <= 24'hff0000;
		12'd1133: rd_data_1 <= 24'hff0000;
		12'd1134: rd_data_1 <= 24'hff0000;
		12'd1135: rd_data_1 <= 24'hff0000;
		12'd1136: rd_data_1 <= 24'h0000ff;
		12'd1137: rd_data_1 <= 24'h0000ff;
		12'd1138: rd_data_1 <= 24'h0000ff;
		12'd1139: rd_data_1 <= 24'h0000ff;
		12'd1140: rd_data_1 <= 24'h0000ff;
		12'd1141: rd_data_1 <= 24'h0000ff;
		12'd1142: rd_data_1 <= 24'h0000ff;
		12'd1143: rd_data_1 <= 24'h0000ff;
		12'd1144: rd_data_1 <= 24'h000000;
		12'd1145: rd_data_1 <= 24'h000000;
		12'd1146: rd_data_1 <= 24'h000000;
		12'd1147: rd_data_1 <= 24'h000000;
		12'd1148: rd_data_1 <= 24'h000000;
		12'd1149: rd_data_1 <= 24'h000000;
		12'd1150: rd_data_1 <= 24'h000000;
		12'd1151: rd_data_1 <= 24'h000000;
		12'd1152: rd_data_1 <= 24'hffffff;
		12'd1153: rd_data_1 <= 24'hffffff;
		12'd1154: rd_data_1 <= 24'hffffff;
		12'd1155: rd_data_1 <= 24'hffffff;
		12'd1156: rd_data_1 <= 24'hffffff;
		12'd1157: rd_data_1 <= 24'hffffff;
		12'd1158: rd_data_1 <= 24'hffffff;
		12'd1159: rd_data_1 <= 24'hffffff;
		12'd1160: rd_data_1 <= 24'hffff00;
		12'd1161: rd_data_1 <= 24'hffff00;
		12'd1162: rd_data_1 <= 24'hffff00;
		12'd1163: rd_data_1 <= 24'hffff00;
		12'd1164: rd_data_1 <= 24'hffff00;
		12'd1165: rd_data_1 <= 24'hffff00;
		12'd1166: rd_data_1 <= 24'hffff00;
		12'd1167: rd_data_1 <= 24'hffff00;
		12'd1168: rd_data_1 <= 24'h00ffff;
		12'd1169: rd_data_1 <= 24'h00ffff;
		12'd1170: rd_data_1 <= 24'h00ffff;
		12'd1171: rd_data_1 <= 24'h00ffff;
		12'd1172: rd_data_1 <= 24'h00ffff;
		12'd1173: rd_data_1 <= 24'h00ffff;
		12'd1174: rd_data_1 <= 24'h00ffff;
		12'd1175: rd_data_1 <= 24'h00ffff;
		12'd1176: rd_data_1 <= 24'h00ff00;
		12'd1177: rd_data_1 <= 24'h00ff00;
		12'd1178: rd_data_1 <= 24'h00ff00;
		12'd1179: rd_data_1 <= 24'h00ff00;
		12'd1180: rd_data_1 <= 24'h00ff00;
		12'd1181: rd_data_1 <= 24'h00ff00;
		12'd1182: rd_data_1 <= 24'h00ff00;
		12'd1183: rd_data_1 <= 24'h00ff00;
		12'd1184: rd_data_1 <= 24'hff00ff;
		12'd1185: rd_data_1 <= 24'hff00ff;
		12'd1186: rd_data_1 <= 24'hff00ff;
		12'd1187: rd_data_1 <= 24'hff00ff;
		12'd1188: rd_data_1 <= 24'hff00ff;
		12'd1189: rd_data_1 <= 24'hff00ff;
		12'd1190: rd_data_1 <= 24'hff00ff;
		12'd1191: rd_data_1 <= 24'hff00ff;
		12'd1192: rd_data_1 <= 24'hff0000;
		12'd1193: rd_data_1 <= 24'hff0000;
		12'd1194: rd_data_1 <= 24'hff0000;
		12'd1195: rd_data_1 <= 24'hff0000;
		12'd1196: rd_data_1 <= 24'hff0000;
		12'd1197: rd_data_1 <= 24'hff0000;
		12'd1198: rd_data_1 <= 24'hff0000;
		12'd1199: rd_data_1 <= 24'hff0000;
		12'd1200: rd_data_1 <= 24'h0000ff;
		12'd1201: rd_data_1 <= 24'h0000ff;
		12'd1202: rd_data_1 <= 24'h0000ff;
		12'd1203: rd_data_1 <= 24'h0000ff;
		12'd1204: rd_data_1 <= 24'h0000ff;
		12'd1205: rd_data_1 <= 24'h0000ff;
		12'd1206: rd_data_1 <= 24'h0000ff;
		12'd1207: rd_data_1 <= 24'h0000ff;
		12'd1208: rd_data_1 <= 24'h000000;
		12'd1209: rd_data_1 <= 24'h000000;
		12'd1210: rd_data_1 <= 24'h000000;
		12'd1211: rd_data_1 <= 24'h000000;
		12'd1212: rd_data_1 <= 24'h000000;
		12'd1213: rd_data_1 <= 24'h000000;
		12'd1214: rd_data_1 <= 24'h000000;
		12'd1215: rd_data_1 <= 24'h000000;
		12'd1216: rd_data_1 <= 24'hffffff;
		12'd1217: rd_data_1 <= 24'hffffff;
		12'd1218: rd_data_1 <= 24'hffffff;
		12'd1219: rd_data_1 <= 24'hffffff;
		12'd1220: rd_data_1 <= 24'hffffff;
		12'd1221: rd_data_1 <= 24'hffffff;
		12'd1222: rd_data_1 <= 24'hffffff;
		12'd1223: rd_data_1 <= 24'hffffff;
		12'd1224: rd_data_1 <= 24'hffff00;
		12'd1225: rd_data_1 <= 24'hffff00;
		12'd1226: rd_data_1 <= 24'hffff00;
		12'd1227: rd_data_1 <= 24'hffff00;
		12'd1228: rd_data_1 <= 24'hffff00;
		12'd1229: rd_data_1 <= 24'hffff00;
		12'd1230: rd_data_1 <= 24'hffff00;
		12'd1231: rd_data_1 <= 24'hffff00;
		12'd1232: rd_data_1 <= 24'h00ffff;
		12'd1233: rd_data_1 <= 24'h00ffff;
		12'd1234: rd_data_1 <= 24'h00ffff;
		12'd1235: rd_data_1 <= 24'h00ffff;
		12'd1236: rd_data_1 <= 24'h00ffff;
		12'd1237: rd_data_1 <= 24'h00ffff;
		12'd1238: rd_data_1 <= 24'h00ffff;
		12'd1239: rd_data_1 <= 24'h00ffff;
		12'd1240: rd_data_1 <= 24'h00ff00;
		12'd1241: rd_data_1 <= 24'h00ff00;
		12'd1242: rd_data_1 <= 24'h00ff00;
		12'd1243: rd_data_1 <= 24'h00ff00;
		12'd1244: rd_data_1 <= 24'h00ff00;
		12'd1245: rd_data_1 <= 24'h00ff00;
		12'd1246: rd_data_1 <= 24'h00ff00;
		12'd1247: rd_data_1 <= 24'h00ff00;
		12'd1248: rd_data_1 <= 24'hff00ff;
		12'd1249: rd_data_1 <= 24'hff00ff;
		12'd1250: rd_data_1 <= 24'hff00ff;
		12'd1251: rd_data_1 <= 24'hff00ff;
		12'd1252: rd_data_1 <= 24'hff00ff;
		12'd1253: rd_data_1 <= 24'hff00ff;
		12'd1254: rd_data_1 <= 24'hff00ff;
		12'd1255: rd_data_1 <= 24'hff00ff;
		12'd1256: rd_data_1 <= 24'hff0000;
		12'd1257: rd_data_1 <= 24'hff0000;
		12'd1258: rd_data_1 <= 24'hff0000;
		12'd1259: rd_data_1 <= 24'hff0000;
		12'd1260: rd_data_1 <= 24'hff0000;
		12'd1261: rd_data_1 <= 24'hff0000;
		12'd1262: rd_data_1 <= 24'hff0000;
		12'd1263: rd_data_1 <= 24'hff0000;
		12'd1264: rd_data_1 <= 24'h0000ff;
		12'd1265: rd_data_1 <= 24'h0000ff;
		12'd1266: rd_data_1 <= 24'h0000ff;
		12'd1267: rd_data_1 <= 24'h0000ff;
		12'd1268: rd_data_1 <= 24'h0000ff;
		12'd1269: rd_data_1 <= 24'h0000ff;
		12'd1270: rd_data_1 <= 24'h0000ff;
		12'd1271: rd_data_1 <= 24'h0000ff;
		12'd1272: rd_data_1 <= 24'h000000;
		12'd1273: rd_data_1 <= 24'h000000;
		12'd1274: rd_data_1 <= 24'h000000;
		12'd1275: rd_data_1 <= 24'h000000;
		12'd1276: rd_data_1 <= 24'h000000;
		12'd1277: rd_data_1 <= 24'h000000;
		12'd1278: rd_data_1 <= 24'h000000;
		12'd1279: rd_data_1 <= 24'h000000;
		12'd1280: rd_data_1 <= 24'hffffff;
		12'd1281: rd_data_1 <= 24'hffffff;
		12'd1282: rd_data_1 <= 24'hffffff;
		12'd1283: rd_data_1 <= 24'hffffff;
		12'd1284: rd_data_1 <= 24'hffffff;
		12'd1285: rd_data_1 <= 24'hffffff;
		12'd1286: rd_data_1 <= 24'hffffff;
		12'd1287: rd_data_1 <= 24'hffffff;
		12'd1288: rd_data_1 <= 24'hffff00;
		12'd1289: rd_data_1 <= 24'hffff00;
		12'd1290: rd_data_1 <= 24'hffff00;
		12'd1291: rd_data_1 <= 24'hffff00;
		12'd1292: rd_data_1 <= 24'hffff00;
		12'd1293: rd_data_1 <= 24'hffff00;
		12'd1294: rd_data_1 <= 24'hffff00;
		12'd1295: rd_data_1 <= 24'hffff00;
		12'd1296: rd_data_1 <= 24'h00ffff;
		12'd1297: rd_data_1 <= 24'h00ffff;
		12'd1298: rd_data_1 <= 24'h00ffff;
		12'd1299: rd_data_1 <= 24'h00ffff;
		12'd1300: rd_data_1 <= 24'h00ffff;
		12'd1301: rd_data_1 <= 24'h00ffff;
		12'd1302: rd_data_1 <= 24'h00ffff;
		12'd1303: rd_data_1 <= 24'h00ffff;
		12'd1304: rd_data_1 <= 24'h00ff00;
		12'd1305: rd_data_1 <= 24'h00ff00;
		12'd1306: rd_data_1 <= 24'h00ff00;
		12'd1307: rd_data_1 <= 24'h00ff00;
		12'd1308: rd_data_1 <= 24'h00ff00;
		12'd1309: rd_data_1 <= 24'h00ff00;
		12'd1310: rd_data_1 <= 24'h00ff00;
		12'd1311: rd_data_1 <= 24'h00ff00;
		12'd1312: rd_data_1 <= 24'hff00ff;
		12'd1313: rd_data_1 <= 24'hff00ff;
		12'd1314: rd_data_1 <= 24'hff00ff;
		12'd1315: rd_data_1 <= 24'hff00ff;
		12'd1316: rd_data_1 <= 24'hff00ff;
		12'd1317: rd_data_1 <= 24'hff00ff;
		12'd1318: rd_data_1 <= 24'hff00ff;
		12'd1319: rd_data_1 <= 24'hff00ff;
		12'd1320: rd_data_1 <= 24'hff0000;
		12'd1321: rd_data_1 <= 24'hff0000;
		12'd1322: rd_data_1 <= 24'hff0000;
		12'd1323: rd_data_1 <= 24'hff0000;
		12'd1324: rd_data_1 <= 24'hff0000;
		12'd1325: rd_data_1 <= 24'hff0000;
		12'd1326: rd_data_1 <= 24'hff0000;
		12'd1327: rd_data_1 <= 24'hff0000;
		12'd1328: rd_data_1 <= 24'h0000ff;
		12'd1329: rd_data_1 <= 24'h0000ff;
		12'd1330: rd_data_1 <= 24'h0000ff;
		12'd1331: rd_data_1 <= 24'h0000ff;
		12'd1332: rd_data_1 <= 24'h0000ff;
		12'd1333: rd_data_1 <= 24'h0000ff;
		12'd1334: rd_data_1 <= 24'h0000ff;
		12'd1335: rd_data_1 <= 24'h0000ff;
		12'd1336: rd_data_1 <= 24'h000000;
		12'd1337: rd_data_1 <= 24'h000000;
		12'd1338: rd_data_1 <= 24'h000000;
		12'd1339: rd_data_1 <= 24'h000000;
		12'd1340: rd_data_1 <= 24'h000000;
		12'd1341: rd_data_1 <= 24'h000000;
		12'd1342: rd_data_1 <= 24'h000000;
		12'd1343: rd_data_1 <= 24'h000000;
		12'd1344: rd_data_1 <= 24'hffffff;
		12'd1345: rd_data_1 <= 24'hffffff;
		12'd1346: rd_data_1 <= 24'hffffff;
		12'd1347: rd_data_1 <= 24'hffffff;
		12'd1348: rd_data_1 <= 24'hffffff;
		12'd1349: rd_data_1 <= 24'hffffff;
		12'd1350: rd_data_1 <= 24'hffffff;
		12'd1351: rd_data_1 <= 24'hffffff;
		12'd1352: rd_data_1 <= 24'hffff00;
		12'd1353: rd_data_1 <= 24'hffff00;
		12'd1354: rd_data_1 <= 24'hffff00;
		12'd1355: rd_data_1 <= 24'hffff00;
		12'd1356: rd_data_1 <= 24'hffff00;
		12'd1357: rd_data_1 <= 24'hffff00;
		12'd1358: rd_data_1 <= 24'hffff00;
		12'd1359: rd_data_1 <= 24'hffff00;
		12'd1360: rd_data_1 <= 24'h00ffff;
		12'd1361: rd_data_1 <= 24'h00ffff;
		12'd1362: rd_data_1 <= 24'h00ffff;
		12'd1363: rd_data_1 <= 24'h00ffff;
		12'd1364: rd_data_1 <= 24'h00ffff;
		12'd1365: rd_data_1 <= 24'h00ffff;
		12'd1366: rd_data_1 <= 24'h00ffff;
		12'd1367: rd_data_1 <= 24'h00ffff;
		12'd1368: rd_data_1 <= 24'h00ff00;
		12'd1369: rd_data_1 <= 24'h00ff00;
		12'd1370: rd_data_1 <= 24'h00ff00;
		12'd1371: rd_data_1 <= 24'h00ff00;
		12'd1372: rd_data_1 <= 24'h00ff00;
		12'd1373: rd_data_1 <= 24'h00ff00;
		12'd1374: rd_data_1 <= 24'h00ff00;
		12'd1375: rd_data_1 <= 24'h00ff00;
		12'd1376: rd_data_1 <= 24'hff00ff;
		12'd1377: rd_data_1 <= 24'hff00ff;
		12'd1378: rd_data_1 <= 24'hff00ff;
		12'd1379: rd_data_1 <= 24'hff00ff;
		12'd1380: rd_data_1 <= 24'hff00ff;
		12'd1381: rd_data_1 <= 24'hff00ff;
		12'd1382: rd_data_1 <= 24'hff00ff;
		12'd1383: rd_data_1 <= 24'hff00ff;
		12'd1384: rd_data_1 <= 24'hff0000;
		12'd1385: rd_data_1 <= 24'hff0000;
		12'd1386: rd_data_1 <= 24'hff0000;
		12'd1387: rd_data_1 <= 24'hff0000;
		12'd1388: rd_data_1 <= 24'hff0000;
		12'd1389: rd_data_1 <= 24'hff0000;
		12'd1390: rd_data_1 <= 24'hff0000;
		12'd1391: rd_data_1 <= 24'hff0000;
		12'd1392: rd_data_1 <= 24'h0000ff;
		12'd1393: rd_data_1 <= 24'h0000ff;
		12'd1394: rd_data_1 <= 24'h0000ff;
		12'd1395: rd_data_1 <= 24'h0000ff;
		12'd1396: rd_data_1 <= 24'h0000ff;
		12'd1397: rd_data_1 <= 24'h0000ff;
		12'd1398: rd_data_1 <= 24'h0000ff;
		12'd1399: rd_data_1 <= 24'h0000ff;
		12'd1400: rd_data_1 <= 24'h000000;
		12'd1401: rd_data_1 <= 24'h000000;
		12'd1402: rd_data_1 <= 24'h000000;
		12'd1403: rd_data_1 <= 24'h000000;
		12'd1404: rd_data_1 <= 24'h000000;
		12'd1405: rd_data_1 <= 24'h000000;
		12'd1406: rd_data_1 <= 24'h000000;
		12'd1407: rd_data_1 <= 24'h000000;
		12'd1408: rd_data_1 <= 24'hffffff;
		12'd1409: rd_data_1 <= 24'hffffff;
		12'd1410: rd_data_1 <= 24'hffffff;
		12'd1411: rd_data_1 <= 24'hffffff;
		12'd1412: rd_data_1 <= 24'hffffff;
		12'd1413: rd_data_1 <= 24'hffffff;
		12'd1414: rd_data_1 <= 24'hffffff;
		12'd1415: rd_data_1 <= 24'hffffff;
		12'd1416: rd_data_1 <= 24'hffff00;
		12'd1417: rd_data_1 <= 24'hffff00;
		12'd1418: rd_data_1 <= 24'hffff00;
		12'd1419: rd_data_1 <= 24'hffff00;
		12'd1420: rd_data_1 <= 24'hffff00;
		12'd1421: rd_data_1 <= 24'hffff00;
		12'd1422: rd_data_1 <= 24'hffff00;
		12'd1423: rd_data_1 <= 24'hffff00;
		12'd1424: rd_data_1 <= 24'h00ffff;
		12'd1425: rd_data_1 <= 24'h00ffff;
		12'd1426: rd_data_1 <= 24'h00ffff;
		12'd1427: rd_data_1 <= 24'h00ffff;
		12'd1428: rd_data_1 <= 24'h00ffff;
		12'd1429: rd_data_1 <= 24'h00ffff;
		12'd1430: rd_data_1 <= 24'h00ffff;
		12'd1431: rd_data_1 <= 24'h00ffff;
		12'd1432: rd_data_1 <= 24'h00ff00;
		12'd1433: rd_data_1 <= 24'h00ff00;
		12'd1434: rd_data_1 <= 24'h00ff00;
		12'd1435: rd_data_1 <= 24'h00ff00;
		12'd1436: rd_data_1 <= 24'h00ff00;
		12'd1437: rd_data_1 <= 24'h00ff00;
		12'd1438: rd_data_1 <= 24'h00ff00;
		12'd1439: rd_data_1 <= 24'h00ff00;
		12'd1440: rd_data_1 <= 24'hff00ff;
		12'd1441: rd_data_1 <= 24'hff00ff;
		12'd1442: rd_data_1 <= 24'hff00ff;
		12'd1443: rd_data_1 <= 24'hff00ff;
		12'd1444: rd_data_1 <= 24'hff00ff;
		12'd1445: rd_data_1 <= 24'hff00ff;
		12'd1446: rd_data_1 <= 24'hff00ff;
		12'd1447: rd_data_1 <= 24'hff00ff;
		12'd1448: rd_data_1 <= 24'hff0000;
		12'd1449: rd_data_1 <= 24'hff0000;
		12'd1450: rd_data_1 <= 24'hff0000;
		12'd1451: rd_data_1 <= 24'hff0000;
		12'd1452: rd_data_1 <= 24'hff0000;
		12'd1453: rd_data_1 <= 24'hff0000;
		12'd1454: rd_data_1 <= 24'hff0000;
		12'd1455: rd_data_1 <= 24'hff0000;
		12'd1456: rd_data_1 <= 24'h0000ff;
		12'd1457: rd_data_1 <= 24'h0000ff;
		12'd1458: rd_data_1 <= 24'h0000ff;
		12'd1459: rd_data_1 <= 24'h0000ff;
		12'd1460: rd_data_1 <= 24'h0000ff;
		12'd1461: rd_data_1 <= 24'h0000ff;
		12'd1462: rd_data_1 <= 24'h0000ff;
		12'd1463: rd_data_1 <= 24'h0000ff;
		12'd1464: rd_data_1 <= 24'h000000;
		12'd1465: rd_data_1 <= 24'h000000;
		12'd1466: rd_data_1 <= 24'h000000;
		12'd1467: rd_data_1 <= 24'h000000;
		12'd1468: rd_data_1 <= 24'h000000;
		12'd1469: rd_data_1 <= 24'h000000;
		12'd1470: rd_data_1 <= 24'h000000;
		12'd1471: rd_data_1 <= 24'h000000;
		12'd1472: rd_data_1 <= 24'hffffff;
		12'd1473: rd_data_1 <= 24'hffffff;
		12'd1474: rd_data_1 <= 24'hffffff;
		12'd1475: rd_data_1 <= 24'hffffff;
		12'd1476: rd_data_1 <= 24'hffffff;
		12'd1477: rd_data_1 <= 24'hffffff;
		12'd1478: rd_data_1 <= 24'hffffff;
		12'd1479: rd_data_1 <= 24'hffffff;
		12'd1480: rd_data_1 <= 24'hffff00;
		12'd1481: rd_data_1 <= 24'hffff00;
		12'd1482: rd_data_1 <= 24'hffff00;
		12'd1483: rd_data_1 <= 24'hffff00;
		12'd1484: rd_data_1 <= 24'hffff00;
		12'd1485: rd_data_1 <= 24'hffff00;
		12'd1486: rd_data_1 <= 24'hffff00;
		12'd1487: rd_data_1 <= 24'hffff00;
		12'd1488: rd_data_1 <= 24'h00ffff;
		12'd1489: rd_data_1 <= 24'h00ffff;
		12'd1490: rd_data_1 <= 24'h00ffff;
		12'd1491: rd_data_1 <= 24'h00ffff;
		12'd1492: rd_data_1 <= 24'h00ffff;
		12'd1493: rd_data_1 <= 24'h00ffff;
		12'd1494: rd_data_1 <= 24'h00ffff;
		12'd1495: rd_data_1 <= 24'h00ffff;
		12'd1496: rd_data_1 <= 24'h00ff00;
		12'd1497: rd_data_1 <= 24'h00ff00;
		12'd1498: rd_data_1 <= 24'h00ff00;
		12'd1499: rd_data_1 <= 24'h00ff00;
		12'd1500: rd_data_1 <= 24'h00ff00;
		12'd1501: rd_data_1 <= 24'h00ff00;
		12'd1502: rd_data_1 <= 24'h00ff00;
		12'd1503: rd_data_1 <= 24'h00ff00;
		12'd1504: rd_data_1 <= 24'hff00ff;
		12'd1505: rd_data_1 <= 24'hff00ff;
		12'd1506: rd_data_1 <= 24'hff00ff;
		12'd1507: rd_data_1 <= 24'hff00ff;
		12'd1508: rd_data_1 <= 24'hff00ff;
		12'd1509: rd_data_1 <= 24'hff00ff;
		12'd1510: rd_data_1 <= 24'hff00ff;
		12'd1511: rd_data_1 <= 24'hff00ff;
		12'd1512: rd_data_1 <= 24'hff0000;
		12'd1513: rd_data_1 <= 24'hff0000;
		12'd1514: rd_data_1 <= 24'hff0000;
		12'd1515: rd_data_1 <= 24'hff0000;
		12'd1516: rd_data_1 <= 24'hff0000;
		12'd1517: rd_data_1 <= 24'hff0000;
		12'd1518: rd_data_1 <= 24'hff0000;
		12'd1519: rd_data_1 <= 24'hff0000;
		12'd1520: rd_data_1 <= 24'h0000ff;
		12'd1521: rd_data_1 <= 24'h0000ff;
		12'd1522: rd_data_1 <= 24'h0000ff;
		12'd1523: rd_data_1 <= 24'h0000ff;
		12'd1524: rd_data_1 <= 24'h0000ff;
		12'd1525: rd_data_1 <= 24'h0000ff;
		12'd1526: rd_data_1 <= 24'h0000ff;
		12'd1527: rd_data_1 <= 24'h0000ff;
		12'd1528: rd_data_1 <= 24'h000000;
		12'd1529: rd_data_1 <= 24'h000000;
		12'd1530: rd_data_1 <= 24'h000000;
		12'd1531: rd_data_1 <= 24'h000000;
		12'd1532: rd_data_1 <= 24'h000000;
		12'd1533: rd_data_1 <= 24'h000000;
		12'd1534: rd_data_1 <= 24'h000000;
		12'd1535: rd_data_1 <= 24'h000000;
		12'd1536: rd_data_1 <= 24'hffffff;
		12'd1537: rd_data_1 <= 24'hffffff;
		12'd1538: rd_data_1 <= 24'hffffff;
		12'd1539: rd_data_1 <= 24'hffffff;
		12'd1540: rd_data_1 <= 24'hffffff;
		12'd1541: rd_data_1 <= 24'hffffff;
		12'd1542: rd_data_1 <= 24'hffffff;
		12'd1543: rd_data_1 <= 24'hffffff;
		12'd1544: rd_data_1 <= 24'hffff00;
		12'd1545: rd_data_1 <= 24'hffff00;
		12'd1546: rd_data_1 <= 24'hffff00;
		12'd1547: rd_data_1 <= 24'hffff00;
		12'd1548: rd_data_1 <= 24'hffff00;
		12'd1549: rd_data_1 <= 24'hffff00;
		12'd1550: rd_data_1 <= 24'hffff00;
		12'd1551: rd_data_1 <= 24'hffff00;
		12'd1552: rd_data_1 <= 24'h00ffff;
		12'd1553: rd_data_1 <= 24'h00ffff;
		12'd1554: rd_data_1 <= 24'h00ffff;
		12'd1555: rd_data_1 <= 24'h00ffff;
		12'd1556: rd_data_1 <= 24'h00ffff;
		12'd1557: rd_data_1 <= 24'h00ffff;
		12'd1558: rd_data_1 <= 24'h00ffff;
		12'd1559: rd_data_1 <= 24'h00ffff;
		12'd1560: rd_data_1 <= 24'h00ff00;
		12'd1561: rd_data_1 <= 24'h00ff00;
		12'd1562: rd_data_1 <= 24'h00ff00;
		12'd1563: rd_data_1 <= 24'h00ff00;
		12'd1564: rd_data_1 <= 24'h00ff00;
		12'd1565: rd_data_1 <= 24'h00ff00;
		12'd1566: rd_data_1 <= 24'h00ff00;
		12'd1567: rd_data_1 <= 24'h00ff00;
		12'd1568: rd_data_1 <= 24'hff00ff;
		12'd1569: rd_data_1 <= 24'hff00ff;
		12'd1570: rd_data_1 <= 24'hff00ff;
		12'd1571: rd_data_1 <= 24'hff00ff;
		12'd1572: rd_data_1 <= 24'hff00ff;
		12'd1573: rd_data_1 <= 24'hff00ff;
		12'd1574: rd_data_1 <= 24'hff00ff;
		12'd1575: rd_data_1 <= 24'hff00ff;
		12'd1576: rd_data_1 <= 24'hff0000;
		12'd1577: rd_data_1 <= 24'hff0000;
		12'd1578: rd_data_1 <= 24'hff0000;
		12'd1579: rd_data_1 <= 24'hff0000;
		12'd1580: rd_data_1 <= 24'hff0000;
		12'd1581: rd_data_1 <= 24'hff0000;
		12'd1582: rd_data_1 <= 24'hff0000;
		12'd1583: rd_data_1 <= 24'hff0000;
		12'd1584: rd_data_1 <= 24'h0000ff;
		12'd1585: rd_data_1 <= 24'h0000ff;
		12'd1586: rd_data_1 <= 24'h0000ff;
		12'd1587: rd_data_1 <= 24'h0000ff;
		12'd1588: rd_data_1 <= 24'h0000ff;
		12'd1589: rd_data_1 <= 24'h0000ff;
		12'd1590: rd_data_1 <= 24'h0000ff;
		12'd1591: rd_data_1 <= 24'h0000ff;
		12'd1592: rd_data_1 <= 24'h000000;
		12'd1593: rd_data_1 <= 24'h000000;
		12'd1594: rd_data_1 <= 24'h000000;
		12'd1595: rd_data_1 <= 24'h000000;
		12'd1596: rd_data_1 <= 24'h000000;
		12'd1597: rd_data_1 <= 24'h000000;
		12'd1598: rd_data_1 <= 24'h000000;
		12'd1599: rd_data_1 <= 24'h000000;
		12'd1600: rd_data_1 <= 24'hffffff;
		12'd1601: rd_data_1 <= 24'hffffff;
		12'd1602: rd_data_1 <= 24'hffffff;
		12'd1603: rd_data_1 <= 24'hffffff;
		12'd1604: rd_data_1 <= 24'hffffff;
		12'd1605: rd_data_1 <= 24'hffffff;
		12'd1606: rd_data_1 <= 24'hffffff;
		12'd1607: rd_data_1 <= 24'hffffff;
		12'd1608: rd_data_1 <= 24'hffff00;
		12'd1609: rd_data_1 <= 24'hffff00;
		12'd1610: rd_data_1 <= 24'hffff00;
		12'd1611: rd_data_1 <= 24'hffff00;
		12'd1612: rd_data_1 <= 24'hffff00;
		12'd1613: rd_data_1 <= 24'hffff00;
		12'd1614: rd_data_1 <= 24'hffff00;
		12'd1615: rd_data_1 <= 24'hffff00;
		12'd1616: rd_data_1 <= 24'h00ffff;
		12'd1617: rd_data_1 <= 24'h00ffff;
		12'd1618: rd_data_1 <= 24'h00ffff;
		12'd1619: rd_data_1 <= 24'h00ffff;
		12'd1620: rd_data_1 <= 24'h00ffff;
		12'd1621: rd_data_1 <= 24'h00ffff;
		12'd1622: rd_data_1 <= 24'h00ffff;
		12'd1623: rd_data_1 <= 24'h00ffff;
		12'd1624: rd_data_1 <= 24'h00ff00;
		12'd1625: rd_data_1 <= 24'h00ff00;
		12'd1626: rd_data_1 <= 24'h00ff00;
		12'd1627: rd_data_1 <= 24'h00ff00;
		12'd1628: rd_data_1 <= 24'h00ff00;
		12'd1629: rd_data_1 <= 24'h00ff00;
		12'd1630: rd_data_1 <= 24'h00ff00;
		12'd1631: rd_data_1 <= 24'h00ff00;
		12'd1632: rd_data_1 <= 24'hff00ff;
		12'd1633: rd_data_1 <= 24'hff00ff;
		12'd1634: rd_data_1 <= 24'hff00ff;
		12'd1635: rd_data_1 <= 24'hff00ff;
		12'd1636: rd_data_1 <= 24'hff00ff;
		12'd1637: rd_data_1 <= 24'hff00ff;
		12'd1638: rd_data_1 <= 24'hff00ff;
		12'd1639: rd_data_1 <= 24'hff00ff;
		12'd1640: rd_data_1 <= 24'hff0000;
		12'd1641: rd_data_1 <= 24'hff0000;
		12'd1642: rd_data_1 <= 24'hff0000;
		12'd1643: rd_data_1 <= 24'hff0000;
		12'd1644: rd_data_1 <= 24'hff0000;
		12'd1645: rd_data_1 <= 24'hff0000;
		12'd1646: rd_data_1 <= 24'hff0000;
		12'd1647: rd_data_1 <= 24'hff0000;
		12'd1648: rd_data_1 <= 24'h0000ff;
		12'd1649: rd_data_1 <= 24'h0000ff;
		12'd1650: rd_data_1 <= 24'h0000ff;
		12'd1651: rd_data_1 <= 24'h0000ff;
		12'd1652: rd_data_1 <= 24'h0000ff;
		12'd1653: rd_data_1 <= 24'h0000ff;
		12'd1654: rd_data_1 <= 24'h0000ff;
		12'd1655: rd_data_1 <= 24'h0000ff;
		12'd1656: rd_data_1 <= 24'h000000;
		12'd1657: rd_data_1 <= 24'h000000;
		12'd1658: rd_data_1 <= 24'h000000;
		12'd1659: rd_data_1 <= 24'h000000;
		12'd1660: rd_data_1 <= 24'h000000;
		12'd1661: rd_data_1 <= 24'h000000;
		12'd1662: rd_data_1 <= 24'h000000;
		12'd1663: rd_data_1 <= 24'h000000;
		12'd1664: rd_data_1 <= 24'hffffff;
		12'd1665: rd_data_1 <= 24'hffffff;
		12'd1666: rd_data_1 <= 24'hffffff;
		12'd1667: rd_data_1 <= 24'hffffff;
		12'd1668: rd_data_1 <= 24'hffffff;
		12'd1669: rd_data_1 <= 24'hffffff;
		12'd1670: rd_data_1 <= 24'hffffff;
		12'd1671: rd_data_1 <= 24'hffffff;
		12'd1672: rd_data_1 <= 24'hffff00;
		12'd1673: rd_data_1 <= 24'hffff00;
		12'd1674: rd_data_1 <= 24'hffff00;
		12'd1675: rd_data_1 <= 24'hffff00;
		12'd1676: rd_data_1 <= 24'hffff00;
		12'd1677: rd_data_1 <= 24'hffff00;
		12'd1678: rd_data_1 <= 24'hffff00;
		12'd1679: rd_data_1 <= 24'hffff00;
		12'd1680: rd_data_1 <= 24'h00ffff;
		12'd1681: rd_data_1 <= 24'h00ffff;
		12'd1682: rd_data_1 <= 24'h00ffff;
		12'd1683: rd_data_1 <= 24'h00ffff;
		12'd1684: rd_data_1 <= 24'h00ffff;
		12'd1685: rd_data_1 <= 24'h00ffff;
		12'd1686: rd_data_1 <= 24'h00ffff;
		12'd1687: rd_data_1 <= 24'h00ffff;
		12'd1688: rd_data_1 <= 24'h00ff00;
		12'd1689: rd_data_1 <= 24'h00ff00;
		12'd1690: rd_data_1 <= 24'h00ff00;
		12'd1691: rd_data_1 <= 24'h00ff00;
		12'd1692: rd_data_1 <= 24'h00ff00;
		12'd1693: rd_data_1 <= 24'h00ff00;
		12'd1694: rd_data_1 <= 24'h00ff00;
		12'd1695: rd_data_1 <= 24'h00ff00;
		12'd1696: rd_data_1 <= 24'hff00ff;
		12'd1697: rd_data_1 <= 24'hff00ff;
		12'd1698: rd_data_1 <= 24'hff00ff;
		12'd1699: rd_data_1 <= 24'hff00ff;
		12'd1700: rd_data_1 <= 24'hff00ff;
		12'd1701: rd_data_1 <= 24'hff00ff;
		12'd1702: rd_data_1 <= 24'hff00ff;
		12'd1703: rd_data_1 <= 24'hff00ff;
		12'd1704: rd_data_1 <= 24'hff0000;
		12'd1705: rd_data_1 <= 24'hff0000;
		12'd1706: rd_data_1 <= 24'hff0000;
		12'd1707: rd_data_1 <= 24'hff0000;
		12'd1708: rd_data_1 <= 24'hff0000;
		12'd1709: rd_data_1 <= 24'hff0000;
		12'd1710: rd_data_1 <= 24'hff0000;
		12'd1711: rd_data_1 <= 24'hff0000;
		12'd1712: rd_data_1 <= 24'h0000ff;
		12'd1713: rd_data_1 <= 24'h0000ff;
		12'd1714: rd_data_1 <= 24'h0000ff;
		12'd1715: rd_data_1 <= 24'h0000ff;
		12'd1716: rd_data_1 <= 24'h0000ff;
		12'd1717: rd_data_1 <= 24'h0000ff;
		12'd1718: rd_data_1 <= 24'h0000ff;
		12'd1719: rd_data_1 <= 24'h0000ff;
		12'd1720: rd_data_1 <= 24'h000000;
		12'd1721: rd_data_1 <= 24'h000000;
		12'd1722: rd_data_1 <= 24'h000000;
		12'd1723: rd_data_1 <= 24'h000000;
		12'd1724: rd_data_1 <= 24'h000000;
		12'd1725: rd_data_1 <= 24'h000000;
		12'd1726: rd_data_1 <= 24'h000000;
		12'd1727: rd_data_1 <= 24'h000000;
		12'd1728: rd_data_1 <= 24'hffffff;
		12'd1729: rd_data_1 <= 24'hffffff;
		12'd1730: rd_data_1 <= 24'hffffff;
		12'd1731: rd_data_1 <= 24'hffffff;
		12'd1732: rd_data_1 <= 24'hffffff;
		12'd1733: rd_data_1 <= 24'hffffff;
		12'd1734: rd_data_1 <= 24'hffffff;
		12'd1735: rd_data_1 <= 24'hffffff;
		12'd1736: rd_data_1 <= 24'hffff00;
		12'd1737: rd_data_1 <= 24'hffff00;
		12'd1738: rd_data_1 <= 24'hffff00;
		12'd1739: rd_data_1 <= 24'hffff00;
		12'd1740: rd_data_1 <= 24'hffff00;
		12'd1741: rd_data_1 <= 24'hffff00;
		12'd1742: rd_data_1 <= 24'hffff00;
		12'd1743: rd_data_1 <= 24'hffff00;
		12'd1744: rd_data_1 <= 24'h00ffff;
		12'd1745: rd_data_1 <= 24'h00ffff;
		12'd1746: rd_data_1 <= 24'h00ffff;
		12'd1747: rd_data_1 <= 24'h00ffff;
		12'd1748: rd_data_1 <= 24'h00ffff;
		12'd1749: rd_data_1 <= 24'h00ffff;
		12'd1750: rd_data_1 <= 24'h00ffff;
		12'd1751: rd_data_1 <= 24'h00ffff;
		12'd1752: rd_data_1 <= 24'h00ff00;
		12'd1753: rd_data_1 <= 24'h00ff00;
		12'd1754: rd_data_1 <= 24'h00ff00;
		12'd1755: rd_data_1 <= 24'h00ff00;
		12'd1756: rd_data_1 <= 24'h00ff00;
		12'd1757: rd_data_1 <= 24'h00ff00;
		12'd1758: rd_data_1 <= 24'h00ff00;
		12'd1759: rd_data_1 <= 24'h00ff00;
		12'd1760: rd_data_1 <= 24'hff00ff;
		12'd1761: rd_data_1 <= 24'hff00ff;
		12'd1762: rd_data_1 <= 24'hff00ff;
		12'd1763: rd_data_1 <= 24'hff00ff;
		12'd1764: rd_data_1 <= 24'hff00ff;
		12'd1765: rd_data_1 <= 24'hff00ff;
		12'd1766: rd_data_1 <= 24'hff00ff;
		12'd1767: rd_data_1 <= 24'hff00ff;
		12'd1768: rd_data_1 <= 24'hff0000;
		12'd1769: rd_data_1 <= 24'hff0000;
		12'd1770: rd_data_1 <= 24'hff0000;
		12'd1771: rd_data_1 <= 24'hff0000;
		12'd1772: rd_data_1 <= 24'hff0000;
		12'd1773: rd_data_1 <= 24'hff0000;
		12'd1774: rd_data_1 <= 24'hff0000;
		12'd1775: rd_data_1 <= 24'hff0000;
		12'd1776: rd_data_1 <= 24'h0000ff;
		12'd1777: rd_data_1 <= 24'h0000ff;
		12'd1778: rd_data_1 <= 24'h0000ff;
		12'd1779: rd_data_1 <= 24'h0000ff;
		12'd1780: rd_data_1 <= 24'h0000ff;
		12'd1781: rd_data_1 <= 24'h0000ff;
		12'd1782: rd_data_1 <= 24'h0000ff;
		12'd1783: rd_data_1 <= 24'h0000ff;
		12'd1784: rd_data_1 <= 24'h000000;
		12'd1785: rd_data_1 <= 24'h000000;
		12'd1786: rd_data_1 <= 24'h000000;
		12'd1787: rd_data_1 <= 24'h000000;
		12'd1788: rd_data_1 <= 24'h000000;
		12'd1789: rd_data_1 <= 24'h000000;
		12'd1790: rd_data_1 <= 24'h000000;
		12'd1791: rd_data_1 <= 24'h000000;
		12'd1792: rd_data_1 <= 24'hffffff;
		12'd1793: rd_data_1 <= 24'hffffff;
		12'd1794: rd_data_1 <= 24'hffffff;
		12'd1795: rd_data_1 <= 24'hffffff;
		12'd1796: rd_data_1 <= 24'hffffff;
		12'd1797: rd_data_1 <= 24'hffffff;
		12'd1798: rd_data_1 <= 24'hffffff;
		12'd1799: rd_data_1 <= 24'hffffff;
		12'd1800: rd_data_1 <= 24'hffff00;
		12'd1801: rd_data_1 <= 24'hffff00;
		12'd1802: rd_data_1 <= 24'hffff00;
		12'd1803: rd_data_1 <= 24'hffff00;
		12'd1804: rd_data_1 <= 24'hffff00;
		12'd1805: rd_data_1 <= 24'hffff00;
		12'd1806: rd_data_1 <= 24'hffff00;
		12'd1807: rd_data_1 <= 24'hffff00;
		12'd1808: rd_data_1 <= 24'h00ffff;
		12'd1809: rd_data_1 <= 24'h00ffff;
		12'd1810: rd_data_1 <= 24'h00ffff;
		12'd1811: rd_data_1 <= 24'h00ffff;
		12'd1812: rd_data_1 <= 24'h00ffff;
		12'd1813: rd_data_1 <= 24'h00ffff;
		12'd1814: rd_data_1 <= 24'h00ffff;
		12'd1815: rd_data_1 <= 24'h00ffff;
		12'd1816: rd_data_1 <= 24'h00ff00;
		12'd1817: rd_data_1 <= 24'h00ff00;
		12'd1818: rd_data_1 <= 24'h00ff00;
		12'd1819: rd_data_1 <= 24'h00ff00;
		12'd1820: rd_data_1 <= 24'h00ff00;
		12'd1821: rd_data_1 <= 24'h00ff00;
		12'd1822: rd_data_1 <= 24'h00ff00;
		12'd1823: rd_data_1 <= 24'h00ff00;
		12'd1824: rd_data_1 <= 24'hff00ff;
		12'd1825: rd_data_1 <= 24'hff00ff;
		12'd1826: rd_data_1 <= 24'hff00ff;
		12'd1827: rd_data_1 <= 24'hff00ff;
		12'd1828: rd_data_1 <= 24'hff00ff;
		12'd1829: rd_data_1 <= 24'hff00ff;
		12'd1830: rd_data_1 <= 24'hff00ff;
		12'd1831: rd_data_1 <= 24'hff00ff;
		12'd1832: rd_data_1 <= 24'hff0000;
		12'd1833: rd_data_1 <= 24'hff0000;
		12'd1834: rd_data_1 <= 24'hff0000;
		12'd1835: rd_data_1 <= 24'hff0000;
		12'd1836: rd_data_1 <= 24'hff0000;
		12'd1837: rd_data_1 <= 24'hff0000;
		12'd1838: rd_data_1 <= 24'hff0000;
		12'd1839: rd_data_1 <= 24'hff0000;
		12'd1840: rd_data_1 <= 24'h0000ff;
		12'd1841: rd_data_1 <= 24'h0000ff;
		12'd1842: rd_data_1 <= 24'h0000ff;
		12'd1843: rd_data_1 <= 24'h0000ff;
		12'd1844: rd_data_1 <= 24'h0000ff;
		12'd1845: rd_data_1 <= 24'h0000ff;
		12'd1846: rd_data_1 <= 24'h0000ff;
		12'd1847: rd_data_1 <= 24'h0000ff;
		12'd1848: rd_data_1 <= 24'h000000;
		12'd1849: rd_data_1 <= 24'h000000;
		12'd1850: rd_data_1 <= 24'h000000;
		12'd1851: rd_data_1 <= 24'h000000;
		12'd1852: rd_data_1 <= 24'h000000;
		12'd1853: rd_data_1 <= 24'h000000;
		12'd1854: rd_data_1 <= 24'h000000;
		12'd1855: rd_data_1 <= 24'h000000;
		12'd1856: rd_data_1 <= 24'hffffff;
		12'd1857: rd_data_1 <= 24'hffffff;
		12'd1858: rd_data_1 <= 24'hffffff;
		12'd1859: rd_data_1 <= 24'hffffff;
		12'd1860: rd_data_1 <= 24'hffffff;
		12'd1861: rd_data_1 <= 24'hffffff;
		12'd1862: rd_data_1 <= 24'hffffff;
		12'd1863: rd_data_1 <= 24'hffffff;
		12'd1864: rd_data_1 <= 24'hffff00;
		12'd1865: rd_data_1 <= 24'hffff00;
		12'd1866: rd_data_1 <= 24'hffff00;
		12'd1867: rd_data_1 <= 24'hffff00;
		12'd1868: rd_data_1 <= 24'hffff00;
		12'd1869: rd_data_1 <= 24'hffff00;
		12'd1870: rd_data_1 <= 24'hffff00;
		12'd1871: rd_data_1 <= 24'hffff00;
		12'd1872: rd_data_1 <= 24'h00ffff;
		12'd1873: rd_data_1 <= 24'h00ffff;
		12'd1874: rd_data_1 <= 24'h00ffff;
		12'd1875: rd_data_1 <= 24'h00ffff;
		12'd1876: rd_data_1 <= 24'h00ffff;
		12'd1877: rd_data_1 <= 24'h00ffff;
		12'd1878: rd_data_1 <= 24'h00ffff;
		12'd1879: rd_data_1 <= 24'h00ffff;
		12'd1880: rd_data_1 <= 24'h00ff00;
		12'd1881: rd_data_1 <= 24'h00ff00;
		12'd1882: rd_data_1 <= 24'h00ff00;
		12'd1883: rd_data_1 <= 24'h00ff00;
		12'd1884: rd_data_1 <= 24'h00ff00;
		12'd1885: rd_data_1 <= 24'h00ff00;
		12'd1886: rd_data_1 <= 24'h00ff00;
		12'd1887: rd_data_1 <= 24'h00ff00;
		12'd1888: rd_data_1 <= 24'hff00ff;
		12'd1889: rd_data_1 <= 24'hff00ff;
		12'd1890: rd_data_1 <= 24'hff00ff;
		12'd1891: rd_data_1 <= 24'hff00ff;
		12'd1892: rd_data_1 <= 24'hff00ff;
		12'd1893: rd_data_1 <= 24'hff00ff;
		12'd1894: rd_data_1 <= 24'hff00ff;
		12'd1895: rd_data_1 <= 24'hff00ff;
		12'd1896: rd_data_1 <= 24'hff0000;
		12'd1897: rd_data_1 <= 24'hff0000;
		12'd1898: rd_data_1 <= 24'hff0000;
		12'd1899: rd_data_1 <= 24'hff0000;
		12'd1900: rd_data_1 <= 24'hff0000;
		12'd1901: rd_data_1 <= 24'hff0000;
		12'd1902: rd_data_1 <= 24'hff0000;
		12'd1903: rd_data_1 <= 24'hff0000;
		12'd1904: rd_data_1 <= 24'h0000ff;
		12'd1905: rd_data_1 <= 24'h0000ff;
		12'd1906: rd_data_1 <= 24'h0000ff;
		12'd1907: rd_data_1 <= 24'h0000ff;
		12'd1908: rd_data_1 <= 24'h0000ff;
		12'd1909: rd_data_1 <= 24'h0000ff;
		12'd1910: rd_data_1 <= 24'h0000ff;
		12'd1911: rd_data_1 <= 24'h0000ff;
		12'd1912: rd_data_1 <= 24'h000000;
		12'd1913: rd_data_1 <= 24'h000000;
		12'd1914: rd_data_1 <= 24'h000000;
		12'd1915: rd_data_1 <= 24'h000000;
		12'd1916: rd_data_1 <= 24'h000000;
		12'd1917: rd_data_1 <= 24'h000000;
		12'd1918: rd_data_1 <= 24'h000000;
		12'd1919: rd_data_1 <= 24'h000000;
		12'd1920: rd_data_1 <= 24'hffffff;
		12'd1921: rd_data_1 <= 24'hffffff;
		12'd1922: rd_data_1 <= 24'hffffff;
		12'd1923: rd_data_1 <= 24'hffffff;
		12'd1924: rd_data_1 <= 24'hffffff;
		12'd1925: rd_data_1 <= 24'hffffff;
		12'd1926: rd_data_1 <= 24'hffffff;
		12'd1927: rd_data_1 <= 24'hffffff;
		12'd1928: rd_data_1 <= 24'hffff00;
		12'd1929: rd_data_1 <= 24'hffff00;
		12'd1930: rd_data_1 <= 24'hffff00;
		12'd1931: rd_data_1 <= 24'hffff00;
		12'd1932: rd_data_1 <= 24'hffff00;
		12'd1933: rd_data_1 <= 24'hffff00;
		12'd1934: rd_data_1 <= 24'hffff00;
		12'd1935: rd_data_1 <= 24'hffff00;
		12'd1936: rd_data_1 <= 24'h00ffff;
		12'd1937: rd_data_1 <= 24'h00ffff;
		12'd1938: rd_data_1 <= 24'h00ffff;
		12'd1939: rd_data_1 <= 24'h00ffff;
		12'd1940: rd_data_1 <= 24'h00ffff;
		12'd1941: rd_data_1 <= 24'h00ffff;
		12'd1942: rd_data_1 <= 24'h00ffff;
		12'd1943: rd_data_1 <= 24'h00ffff;
		12'd1944: rd_data_1 <= 24'h00ff00;
		12'd1945: rd_data_1 <= 24'h00ff00;
		12'd1946: rd_data_1 <= 24'h00ff00;
		12'd1947: rd_data_1 <= 24'h00ff00;
		12'd1948: rd_data_1 <= 24'h00ff00;
		12'd1949: rd_data_1 <= 24'h00ff00;
		12'd1950: rd_data_1 <= 24'h00ff00;
		12'd1951: rd_data_1 <= 24'h00ff00;
		12'd1952: rd_data_1 <= 24'hff00ff;
		12'd1953: rd_data_1 <= 24'hff00ff;
		12'd1954: rd_data_1 <= 24'hff00ff;
		12'd1955: rd_data_1 <= 24'hff00ff;
		12'd1956: rd_data_1 <= 24'hff00ff;
		12'd1957: rd_data_1 <= 24'hff00ff;
		12'd1958: rd_data_1 <= 24'hff00ff;
		12'd1959: rd_data_1 <= 24'hff00ff;
		12'd1960: rd_data_1 <= 24'hff0000;
		12'd1961: rd_data_1 <= 24'hff0000;
		12'd1962: rd_data_1 <= 24'hff0000;
		12'd1963: rd_data_1 <= 24'hff0000;
		12'd1964: rd_data_1 <= 24'hff0000;
		12'd1965: rd_data_1 <= 24'hff0000;
		12'd1966: rd_data_1 <= 24'hff0000;
		12'd1967: rd_data_1 <= 24'hff0000;
		12'd1968: rd_data_1 <= 24'h0000ff;
		12'd1969: rd_data_1 <= 24'h0000ff;
		12'd1970: rd_data_1 <= 24'h0000ff;
		12'd1971: rd_data_1 <= 24'h0000ff;
		12'd1972: rd_data_1 <= 24'h0000ff;
		12'd1973: rd_data_1 <= 24'h0000ff;
		12'd1974: rd_data_1 <= 24'h0000ff;
		12'd1975: rd_data_1 <= 24'h0000ff;
		12'd1976: rd_data_1 <= 24'h000000;
		12'd1977: rd_data_1 <= 24'h000000;
		12'd1978: rd_data_1 <= 24'h000000;
		12'd1979: rd_data_1 <= 24'h000000;
		12'd1980: rd_data_1 <= 24'h000000;
		12'd1981: rd_data_1 <= 24'h000000;
		12'd1982: rd_data_1 <= 24'h000000;
		12'd1983: rd_data_1 <= 24'h000000;
		12'd1984: rd_data_1 <= 24'hffffff;
		12'd1985: rd_data_1 <= 24'hffffff;
		12'd1986: rd_data_1 <= 24'hffffff;
		12'd1987: rd_data_1 <= 24'hffffff;
		12'd1988: rd_data_1 <= 24'hffffff;
		12'd1989: rd_data_1 <= 24'hffffff;
		12'd1990: rd_data_1 <= 24'hffffff;
		12'd1991: rd_data_1 <= 24'hffffff;
		12'd1992: rd_data_1 <= 24'hffff00;
		12'd1993: rd_data_1 <= 24'hffff00;
		12'd1994: rd_data_1 <= 24'hffff00;
		12'd1995: rd_data_1 <= 24'hffff00;
		12'd1996: rd_data_1 <= 24'hffff00;
		12'd1997: rd_data_1 <= 24'hffff00;
		12'd1998: rd_data_1 <= 24'hffff00;
		12'd1999: rd_data_1 <= 24'hffff00;
		12'd2000: rd_data_1 <= 24'h00ffff;
		12'd2001: rd_data_1 <= 24'h00ffff;
		12'd2002: rd_data_1 <= 24'h00ffff;
		12'd2003: rd_data_1 <= 24'h00ffff;
		12'd2004: rd_data_1 <= 24'h00ffff;
		12'd2005: rd_data_1 <= 24'h00ffff;
		12'd2006: rd_data_1 <= 24'h00ffff;
		12'd2007: rd_data_1 <= 24'h00ffff;
		12'd2008: rd_data_1 <= 24'h00ff00;
		12'd2009: rd_data_1 <= 24'h00ff00;
		12'd2010: rd_data_1 <= 24'h00ff00;
		12'd2011: rd_data_1 <= 24'h00ff00;
		12'd2012: rd_data_1 <= 24'h00ff00;
		12'd2013: rd_data_1 <= 24'h00ff00;
		12'd2014: rd_data_1 <= 24'h00ff00;
		12'd2015: rd_data_1 <= 24'h00ff00;
		12'd2016: rd_data_1 <= 24'hff00ff;
		12'd2017: rd_data_1 <= 24'hff00ff;
		12'd2018: rd_data_1 <= 24'hff00ff;
		12'd2019: rd_data_1 <= 24'hff00ff;
		12'd2020: rd_data_1 <= 24'hff00ff;
		12'd2021: rd_data_1 <= 24'hff00ff;
		12'd2022: rd_data_1 <= 24'hff00ff;
		12'd2023: rd_data_1 <= 24'hff00ff;
		12'd2024: rd_data_1 <= 24'hff0000;
		12'd2025: rd_data_1 <= 24'hff0000;
		12'd2026: rd_data_1 <= 24'hff0000;
		12'd2027: rd_data_1 <= 24'hff0000;
		12'd2028: rd_data_1 <= 24'hff0000;
		12'd2029: rd_data_1 <= 24'hff0000;
		12'd2030: rd_data_1 <= 24'hff0000;
		12'd2031: rd_data_1 <= 24'hff0000;
		12'd2032: rd_data_1 <= 24'h0000ff;
		12'd2033: rd_data_1 <= 24'h0000ff;
		12'd2034: rd_data_1 <= 24'h0000ff;
		12'd2035: rd_data_1 <= 24'h0000ff;
		12'd2036: rd_data_1 <= 24'h0000ff;
		12'd2037: rd_data_1 <= 24'h0000ff;
		12'd2038: rd_data_1 <= 24'h0000ff;
		12'd2039: rd_data_1 <= 24'h0000ff;
		12'd2040: rd_data_1 <= 24'h000000;
		12'd2041: rd_data_1 <= 24'h000000;
		12'd2042: rd_data_1 <= 24'h000000;
		12'd2043: rd_data_1 <= 24'h000000;
		12'd2044: rd_data_1 <= 24'h000000;
		12'd2045: rd_data_1 <= 24'h000000;
		12'd2046: rd_data_1 <= 24'h000000;
		12'd2047: rd_data_1 <= 24'h000000;

        endcase
    end    
        assign o_rd_data[0][2] = rd_data_0[3*bpp_p-1-:8];
        assign o_rd_data[0][1] = rd_data_0[2*bpp_p-1-:8];
        assign o_rd_data[0][0] = rd_data_0[bpp_p-1-:8];

        assign o_rd_data[1][2] = rd_data_1[3*bpp_p-1-:8];
        assign o_rd_data[1][1] = rd_data_1[2*bpp_p-1-:8];
        assign o_rd_data[1][0] = rd_data_1[bpp_p-1-:8];
endmodule