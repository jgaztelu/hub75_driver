module bulbasaur_rom #(
	parameter hpixel_p = 65,
    parameter vpixel_p = 65,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

// Clock and reset
        input logic clk,
        input logic rst_n,

        /* Pixel read interface */
        input logic [addr_width_p-1:0] i_rd_addr,
        output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
        );

localparam [frame_size_p-1:0][3*bpp_p-1:0] bulbasaur_rom_buf = {
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h810081,
24'h810081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f017c,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f017c,
24'h7f017c,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7d0081,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h81007e,
24'h7f017c,
24'h7f017c,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f0081,
24'h7f0083,
24'h810081,
24'h810081,
24'h7f0081,
24'h7d007f,
24'h7d017e,
24'h7d007d,
24'h830183,
24'h810083,
24'h81007f,
24'h7f007e,
24'h7f007e,
24'h7d017e,
24'h7d017e,
24'h7b017e,
24'h7b017e,
24'h79027c,
24'h750579,
24'h77047b,
24'h7b007f,
24'h7f0081,
24'h81007f,
24'h81007e,
24'h7f017c,
24'h7f017c,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f017c,
24'h7f0477,
24'h7d0379,
24'h7d0083,
24'h7d0083,
24'h7d027c,
24'h7d027c,
24'h7d0084,
24'h810087,
24'h870086,
24'h850084,
24'h7f0083,
24'h7b007f,
24'h800a82,
24'h760077,
24'h88008a,
24'h89008b,
24'h8c0889,
24'h850480,
24'h7e037d,
24'h7a017b,
24'h720078,
24'h71017a,
24'h740880,
24'h670474,
24'h6a1673,
24'h63096c,
24'h72027d,
24'h78007e,
24'h85007e,
24'h85017b,
24'h81027b,
24'h7f017c,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f0379,
24'h7f027b,
24'h7f0084,
24'h7f0084,
24'h7f027b,
24'h7f027b,
24'h7f0083,
24'h830086,
24'h870086,
24'h870084,
24'h810081,
24'h7b007b,
24'h740075,
24'h750076,
24'h830383,
24'h7d007a,
24'h7a0972,
24'h6a0260,
24'h690563,
24'h751673,
24'h630b67,
24'h6d1a75,
24'h65156f,
24'h561562,
24'h4c2556,
24'h62386a,
24'h5e1265,
24'h610065,
24'h7a0573,
24'h7f0477,
24'h7d037b,
24'h7d027c,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h81007e,
24'h81007e,
24'h81007f,
24'h81007f,
24'h81007f,
24'h81007f,
24'h81007e,
24'h81007f,
24'h830084,
24'h830083,
24'h83017b,
24'h840479,
24'h85007c,
24'h85007f,
24'h850083,
24'h850081,
24'h87007c,
24'h87027f,
24'h860484,
24'h7e067e,
24'h6d0568,
24'h6d1563,
24'h692259,
24'h5d214b,
24'h562048,
24'h55234b,
24'h481d44,
24'h4e284e,
24'h442046,
24'h564759,
24'h394f3d,
24'h8da48e,
24'h12090f,
24'h2c0029,
24'h5c0f60,
24'h6f0974,
24'h750579,
24'h79027c,
24'h7d017e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h81007e,
24'h81007e,
24'h81007f,
24'h81007f,
24'h81007f,
24'h81007f,
24'h81007e,
24'h81007f,
24'h83007f,
24'h83007f,
24'h810078,
24'h84037a,
24'h85017b,
24'h83017c,
24'h81007f,
24'h81007f,
24'h83017b,
24'h7f0576,
24'h780c75,
24'h640f64,
24'h582052,
24'h816078,
24'h857174,
24'h8a7e79,
24'h766e69,
24'h514f48,
24'h4d524a,
24'h464f47,
24'h455148,
24'h8ba88f,
24'h4b8651,
24'h518b52,
24'h415c3a,
24'h766a71,
24'h460c4a,
24'h660b6e,
24'h730375,
24'h7d027c,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7a0076,
24'h870c80,
24'h77006f,
24'h80047a,
24'h7a0078,
24'h810380,
24'h750072,
24'h81047f,
24'h840786,
24'h810988,
24'h7a0881,
24'h670b6c,
24'h592357,
24'h796977,
24'h647a69,
24'ha3cca5,
24'habd1a4,
24'ha6cd9e,
24'ha0cb9b,
24'h9ece9e,
24'ha0d8a6,
24'h7db986,
24'h70af7c,
24'h77ba84,
24'h45894e,
24'h7cb57e,
24'h3f613a,
24'h6f6f6a,
24'h2d002d,
24'h731771,
24'h7a0071,
24'h8f0884,
24'h82017f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d0477,
24'h831774,
24'h7c1664,
24'h710d58,
24'h7c1469,
24'h75066f,
24'h7a0a79,
24'h790977,
24'h7e0e7b,
24'h7b0d7a,
24'h751077,
24'h67126d,
24'h511954,
24'h7f6f76,
24'hbaceaf,
24'haadca4,
24'h9fdd98,
24'ha4de97,
24'ha1db94,
24'h9bda93,
24'h9ade95,
24'h90d88f,
24'h9ae79d,
24'h3b8d42,
24'h43924a,
24'h80c781,
24'h82be7f,
24'h5a8353,
24'h4d5748,
24'h21001e,
24'h60105c,
24'h7f0574,
24'h89007e,
24'h840081,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h790a6e,
24'h6a1a44,
24'h6c2939,
24'h763542,
24'h6d2643,
24'h721f5e,
24'h6b1361,
24'h6e1765,
24'h660e5c,
24'h64105b,
24'h57114d,
24'h5f3351,
24'h857172,
24'hc2c7ab,
24'hb5ca99,
24'hb3d390,
24'hb5dc91,
24'hb2da92,
24'h2b550f,
24'h023100,
24'h4d8139,
24'h559047,
24'h4d8d43,
24'h9ddf95,
24'h7dc373,
24'h74ba64,
24'h7bba69,
24'h598a50,
24'h435a3e,
24'h1b0a14,
24'h5c2158,
24'h7a0c79,
24'h88058a,
24'h800082,
24'h800181,
24'h820082,
24'h820082,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h750e67,
24'hab717a,
24'hf2d2b1,
24'hedd1aa,
24'h6a4931,
24'h60343d,
24'h62304a,
24'h86526b,
24'h88556b,
24'h805164,
24'h7d595d,
24'h6f6448,
24'h69703f,
24'h6a7d3d,
24'h587227,
24'h5c7425,
24'h375202,
24'h3c5b0d,
24'hc0e298,
24'hadce8d,
24'h062d00,
24'h9ccc89,
24'h9ed78e,
24'h98d98c,
24'h98de8a,
24'h82c969,
24'h78bb61,
24'h7fb972,
24'h3d6435,
24'h747d67,
24'h290b20,
24'h601162,
24'h700074,
24'h7e0181,
24'h820082,
24'h820082,
24'h820082,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d007f,
24'h7d0081,
24'h711064,
24'h99776a,
24'he5e5a1,
24'hd0de8c,
24'hd7e797,
24'h6b7339,
24'h656737,
24'hd8d2a1,
24'hdcd8a2,
24'hd8d89c,
24'hd4db98,
24'hd8e996,
24'hb9d373,
24'hb2d069,
24'hb4d26b,
24'h3d5800,
24'hd0ec93,
24'hcaed93,
24'hc7e79b,
24'hb4c89a,
24'h0b2000,
24'hadd49d,
24'h9ed591,
24'h92dd8d,
24'h8ddd84,
24'h79c368,
24'h7abf64,
24'h7bc06e,
24'h387329,
24'h5e8548,
24'h757d60,
24'h290322,
24'h6a1b6a,
24'h7b037b,
24'h860085,
24'h840084,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d0081,
24'h6f1261,
24'h998268,
24'hd0e28b,
24'h7ea139,
24'hbde67b,
24'hc4e88c,
24'hcdeb92,
24'hcee284,
24'hd1e483,
24'h7e9536,
24'h7f9938,
24'h7e9b32,
24'hd3f282,
24'hb6d95d,
24'hb0d259,
24'hc2de75,
24'hc6e381,
24'hc5ea84,
24'habcb74,
24'hb2c48f,
24'h0d2000,
24'hb7d7a6,
24'h9ed192,
24'h96e393,
24'h93e88f,
24'h78c36e,
24'h7ec36f,
24'h76c06b,
24'h408531,
24'h316816,
24'h719057,
24'h221b13,
24'h521e4d,
24'h750873,
24'h840084,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7b017e,
24'h7b007f,
24'h7b007f,
24'h7b007f,
24'h7b027c,
24'h6d165b,
24'h998561,
24'h667a1e,
24'hc7ea82,
24'hcbf38b,
24'hc7eb8c,
24'hc6e686,
24'hd2ec7f,
24'h8aa134,
24'h899f43,
24'h7d943c,
24'h859d42,
24'hceeb82,
24'hcff473,
24'hb4d956,
24'hbbda69,
24'hb2d166,
24'hb9dd6c,
24'hadcf65,
24'hacc56d,
24'h7a924c,
24'h092500,
24'ha1cf98,
24'h9ae294,
24'h92e38d,
24'h7bc276,
24'h80c47b,
24'h75bb6b,
24'h4f913f,
24'h336d18,
24'h6a914d,
24'h697656,
24'h26091b,
24'h691067,
24'h7c037d,
24'h800181,
24'h820082,
24'h820082,
24'h820082,
24'h820082,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7b027c,
24'h7b017e,
24'h7b0081,
24'h7b017e,
24'h7b0577,
24'h6d1954,
24'h837048,
24'hcde281,
24'hc4e77d,
24'hb7df77,
24'hc7ea8e,
24'hcbea8c,
24'h8aa338,
24'h7e9529,
24'h839a3c,
24'h768e33,
24'hc6de83,
24'hd4f089,
24'hd3f778,
24'hbde162,
24'ha9c65b,
24'hb5d06c,
24'hb6d867,
24'hb5d562,
24'hb8d466,
24'h768f37,
24'h061f00,
24'hadd5a3,
24'h98db8e,
24'h80cb79,
24'h79c07a,
24'h7fc480,
24'h7ac072,
24'h4d903e,
24'h548e3c,
24'h34641a,
24'h62844d,
24'h16120a,
24'h5d185c,
24'h740877,
24'h7b027c,
24'h800181,
24'h830083,
24'h830083,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d027c,
24'h7b037b,
24'h7b027c,
24'h79007f,
24'h7a007d,
24'h7c0972,
24'h69194a,
24'h79683d,
24'hcae07f,
24'hc8ee7f,
24'hcbf489,
24'hccef95,
24'hbeda86,
24'h84973e,
24'h859739,
24'h87a03a,
24'hd1ed84,
24'hceeb82,
24'hd4f286,
24'hd4f383,
24'hbbd76e,
24'h879d49,
24'h798e3d,
24'hb3cb6a,
24'hb3cc5f,
24'hc1da66,
24'h859d3a,
24'h0c2100,
24'hb4d4a6,
24'h80bb72,
24'h78c171,
24'h7ac17c,
24'h7bc27d,
24'h599d4e,
24'h539440,
24'h528d3d,
24'h366e20,
24'h568f44,
24'h6f8664,
24'h2f002f,
24'h690d6e,
24'h750677,
24'h7c007c,
24'h830083,
24'h830083,
24'h7f007f,
24'h7d017e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d027c,
24'h7b037b,
24'h7b027c,
24'h75007b,
24'h7d047f,
24'h790968,
24'h914170,
24'h5b4530,
24'hd0df98,
24'haacb69,
24'hbee67e,
24'hc0e387,
24'hc8e38c,
24'hd1e28f,
24'hd7e690,
24'hc6df79,
24'hd3f184,
24'hcbe97b,
24'hb6d06e,
24'hd2e49a,
24'h6a7541,
24'hd2d5b7,
24'hd5d8b3,
24'h4c5610,
24'hbfcf71,
24'h8d9f33,
24'h899c3b,
24'h7a8851,
24'h0b2600,
24'h82b771,
24'h79bf70,
24'h72bd73,
24'h428f40,
24'h549b42,
24'h4c8b34,
24'h549042,
24'h2d6b1f,
24'h539b46,
24'h547d4d,
24'h230527,
24'h611267,
24'h720675,
24'h7c007a,
24'h840083,
24'h840083,
24'h7c007d,
24'h7a017b,
24'h7d017e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d027c,
24'h7d0379,
24'h7d037b,
24'h7c0084,
24'h7c047c,
24'h790b64,
24'h712059,
24'h745169,
24'h838270,
24'hc1d993,
24'hb0d675,
24'hcdf18e,
24'hcae686,
24'hd4e48d,
24'h8c9943,
24'h809836,
24'hc9e47e,
24'hb0cc65,
24'hd2e39c,
24'h5f5951,
24'h665273,
24'h41295d,
24'hffefff,
24'hdfd7bb,
24'h525510,
24'h8d933e,
24'h7a8332,
24'h808a52,
24'h061c00,
24'h2d5d1a,
24'h599a4c,
24'h43923d,
24'h4fa144,
24'h4e9835,
24'h498b2e,
24'h5a954a,
24'h2a6b23,
24'h3e913d,
24'h528854,
24'h190a21,
24'h5b1563,
24'h700871,
24'h7c007a,
24'h860083,
24'h840083,
24'h7c007d,
24'h7a017b,
24'h7d017e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h7d017e,
24'h7d027c,
24'h7d037b,
24'h7d027c,
24'h76007c,
24'h760673,
24'h701859,
24'h682956,
24'h6b477b,
24'h81788c,
24'hcadea9,
24'hafd173,
24'hc8ec82,
24'hcfeb85,
24'h86943b,
24'h7e8b35,
24'h789132,
24'hcbe886,
24'hb1cb6b,
24'hd5dcab,
24'h6b5679,
24'h623d97,
24'h3c1484,
24'hffe2ff,
24'hfffdfd,
24'h534c16,
24'h959649,
24'h8a8f3c,
24'h7f8544,
24'h1b2b00,
24'h32520f,
24'h5d9142,
24'h4b923a,
24'h499436,
24'h4b8f30,
24'h57973f,
24'h347127,
24'h478b42,
24'h449645,
24'h4f8152,
24'h1f0726,
24'h611366,
24'h720773,
24'h7c007a,
24'h840083,
24'h840083,
24'h7c007d,
24'h7a017b,
24'h7d017e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f017c,
24'h7f027b,
24'h7f017c,
24'h7d017e,
24'h79007b,
24'h6d0c67,
24'h80546b,
24'hdbc3d3,
24'h694d8c,
24'hfcedff,
24'h7a895e,
24'hc4e385,
24'hd2f286,
24'hd7f085,
24'h8d9842,
24'h8a9642,
24'hc4e47f,
24'hcef08b,
24'hcee28c,
24'h8b8869,
24'h674785,
24'hffd4ff,
24'h320695,
24'h391783,
24'hfff7ff,
24'he3daab,
24'h8e9137,
24'h9aa23f,
24'h8a9140,
24'h49510c,
24'h7d8741,
24'h3e580b,
24'h5c8f37,
24'h57923b,
24'h528a3c,
24'h629a51,
24'h2b671b,
24'h4a8a40,
24'h50964d,
24'h5c785c,
24'h350037,
24'h6f0471,
24'h820d82,
24'h780079,
24'h81007f,
24'h81007f,
24'h7d017e,
24'h7d027c,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f027b,
24'h7f027b,
24'h7f017c,
24'h7f007e,
24'h7c017b,
24'h660a5d,
24'h755a5a,
24'hfffef5,
24'h39245b,
24'hfcedff,
24'h7a8b59,
24'hb8d871,
24'hceee7c,
24'hd8f081,
24'hd4e184,
24'hd5e587,
24'hd4f68a,
24'hc7e87f,
24'hbcce77,
24'h858361,
24'h43295d,
24'hffe0ff,
24'h9779f2,
24'h8d75cf,
24'hfff4ff,
24'he8deb0,
24'h94963f,
24'h89932d,
24'h929a40,
24'h767a2a,
24'h94934b,
24'h878e44,
24'h395300,
24'h709542,
24'h648a42,
24'h3c6821,
24'h4d893b,
24'h529149,
24'h4f804d,
24'h101010,
24'h610f61,
24'h7f047f,
24'h800781,
24'h7e037d,
24'h7f007e,
24'h7f007e,
24'h7d027c,
24'h7d027c,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h81017c,
24'h81027b,
24'h7f027b,
24'h7f027b,
24'h78007b,
24'h76186b,
24'h815e5a,
24'hc0b8a2,
24'h3c2d4d,
24'h332e3d,
24'h788f43,
24'hb4d85e,
24'hb7d75c,
24'hb7d25a,
24'hc1d867,
24'hbed463,
24'hb3d057,
24'hb6d25e,
24'hb8cd68,
24'h888e52,
24'h3c3437,
24'h3b325a,
24'h8889b6,
24'h8a8ca7,
24'hd8d0bf,
24'h8f8756,
24'h99984f,
24'h949841,
24'h939a3b,
24'h8f943b,
24'h8d8c44,
24'h908f49,
24'h909244,
24'h505704,
24'h495705,
24'h6e8f3c,
24'h62a14b,
24'h53904f,
24'h5d705f,
24'h25072a,
24'h741774,
24'h810580,
24'h7f047f,
24'h820681,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h81007f,
24'h83007e,
24'h83017c,
24'h7f0379,
24'h7f027b,
24'h810282,
24'h78136c,
24'h633339,
24'h281600,
24'hb6a9b0,
24'haeaca5,
24'hb8c58a,
24'hb7d071,
24'hb7d364,
24'hbbd861,
24'hb7d15d,
24'hbad261,
24'hbad35f,
24'hbfd768,
24'hbcd26f,
24'hb9c881,
24'hadb49a,
24'hafb7af,
24'h97a99d,
24'ha0af98,
24'h83825c,
24'h968f5a,
24'h54520e,
24'h8b8d3d,
24'h8d9337,
24'h8f943b,
24'h97984d,
24'h97934d,
24'h968f47,
24'h9c954b,
24'h969848,
24'h455909,
24'h5a9041,
24'h5e8759,
24'h190819,
24'h642266,
24'h6c046e,
24'h7e037d,
24'h820681,
24'h7e037d,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h81007f,
24'h85007f,
24'h85007e,
24'h7f0379,
24'h7d037b,
24'h7c007c,
24'h760a6b,
24'h6b2749,
24'h9b7771,
24'h201300,
24'h413b2a,
24'hbcb1b1,
24'hc2c0ac,
24'h839648,
24'hb6d368,
24'hc2dc76,
24'h667f1b,
24'hadc662,
24'hbbd376,
24'hadc374,
24'habc082,
24'ha4b58b,
24'hb5c7a0,
24'h596c39,
24'h3a480f,
24'h202100,
24'h211d00,
24'h8e8e45,
24'h898b3b,
24'h727424,
24'h929444,
24'h8e9040,
24'h878940,
24'h4f4f11,
24'h515015,
24'h92914f,
24'h838c48,
24'h335015,
24'h171b08,
24'h612257,
24'h6f076a,
24'h790479,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h870083,
24'h870081,
24'h7f017c,
24'h7d037b,
24'h80027f,
24'h7e0a76,
24'h630a4f,
24'h652a46,
24'h947b6f,
24'hffffef,
24'h3c2938,
24'h403337,
24'hb4bc8f,
24'hb6c58c,
24'hb4bb98,
24'hb7bba2,
24'hadb49a,
24'h656d57,
24'h3e473a,
24'h121e10,
24'h091702,
24'h0e1b00,
24'hffffd1,
24'h6a7028,
24'h8e8e50,
24'h8e8b51,
24'h93914d,
24'h909047,
24'h57590b,
24'h8b8d3d,
24'h949947,
24'h8e9347,
24'h52561a,
24'h4e5218,
24'h525313,
24'h909453,
24'h79854f,
24'h4a3d2f,
24'h6b215a,
24'h6e0165,
24'h7b0479,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h830081,
24'h890084,
24'h870084,
24'h7f0081,
24'h7b017e,
24'h7c0076,
24'h85097f,
24'h7a0a79,
24'h691264,
24'h5a2c4a,
24'h927c79,
24'h8c806d,
24'h686450,
24'h3a3630,
24'h362845,
24'h3c1e70,
24'h421f8b,
24'h2d1179,
24'h30197f,
24'h2b1a7c,
24'h2b216e,
24'h332d53,
24'h433c37,
24'h796f3c,
24'h938941,
24'h918a47,
24'h989253,
24'h978e59,
24'h4f4b0e,
24'h8e913e,
24'h91983e,
24'h89913d,
24'h979f52,
24'h879048,
24'h4e5610,
24'h4c5208,
24'h888b44,
24'h8c8f4f,
24'h8e8060,
24'h64324d,
24'h67155e,
24'h750873,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h870084,
24'h850084,
24'h7d0083,
24'h7d007f,
24'h790072,
24'h7c0078,
24'h7c0084,
24'h6f0377,
24'h6c226a,
24'h360524,
24'h33130d,
24'h927e6f,
24'h817176,
24'h604e76,
24'h33126c,
24'h633fb2,
24'h926fe4,
24'h8d72e4,
24'h816dd9,
24'h8277c8,
24'h605a82,
24'h807875,
24'h918454,
24'h998a44,
24'ha49954,
24'h2b2200,
24'h342900,
24'h8e8849,
24'h898f38,
24'h919c3f,
24'h858e3d,
24'h869043,
24'h6e7829,
24'h889344,
24'h8a9246,
24'h8c9147,
24'h94934c,
24'h918454,
24'h583834,
24'h561945,
24'h730b6e,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h810081,
24'h810081,
24'h7d0081,
24'h7d007f,
24'h80007b,
24'h80007d,
24'h7e0081,
24'h7a0080,
24'h78097b,
24'h6e0e66,
24'h6c1a50,
24'h370011,
24'h1c0c00,
24'h86866b,
24'h7c7c6e,
24'h7d7978,
24'h807280,
24'h7c7183,
24'h7c7c8a,
24'h7c8487,
24'h758373,
24'h7e8a66,
24'h282700,
24'h2c2500,
24'h312300,
24'h968a4a,
24'h928c3f,
24'h868831,
24'h70771f,
24'h838b36,
24'h848d43,
24'h495409,
24'h86963f,
24'h87943e,
24'h8a8e45,
24'h50500c,
24'h8b8842,
24'h91844b,
24'h998064,
24'h3e071c,
24'h730e67,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7f007f,
24'h7e007d,
24'h80007d,
24'h7e0081,
24'h7e0083,
24'h73007a,
24'h7e047c,
24'h760863,
24'h762c53,
24'h948261,
24'h1d2a00,
24'h1d3000,
24'h111f00,
24'h222200,
24'h262600,
24'h161f00,
24'h0d2000,
24'h0d2500,
24'h0c1f00,
24'h858c48,
24'h92904a,
24'h928a43,
24'h958d3f,
24'h918f35,
24'h909234,
24'h4e5400,
24'h888d41,
24'h8a8e4e,
24'h282f00,
24'h859136,
24'h909a40,
24'h575811,
24'h575415,
24'h56510f,
24'h887d44,
24'h9c8a62,
24'h400f17,
24'h730f66,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7e007d,
24'h7e007d,
24'h7e0081,
24'h7e0083,
24'h7e0084,
24'h750074,
24'h7e0c73,
24'hab5e8c,
24'hcabc8e,
24'hb0c264,
24'hb6cc6b,
24'h86963f,
24'h4d510e,
24'h888c52,
24'h859355,
24'h7f924d,
24'h869b48,
24'h7d8c37,
24'h8f934a,
24'h4c4e00,
24'hced36b,
24'hcace62,
24'h969937,
24'h8e9039,
24'h8d8e41,
24'h535311,
24'h1a1600,
24'h89864b,
24'h959b3f,
24'h868a2c,
24'h57530f,
24'h504810,
24'h524c12,
24'h8e8653,
24'h8b815c,
24'h2a010a,
24'h710f66,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7e007d,
24'h7e007d,
24'h7e0081,
24'h7e0081,
24'h86098a,
24'h780079,
24'h7d077a,
24'h6c1c54,
24'h7e6d40,
24'h859634,
24'hb8ce66,
24'hb6c969,
24'h848a3c,
24'h4e4f0d,
24'h252f00,
24'h7b8447,
24'h89884d,
24'h888545,
24'h4c4d06,
24'h919742,
24'h939e33,
24'hc3cd5f,
24'hccd26f,
24'h8d8f38,
24'h8d8c44,
24'h575119,
24'h291b00,
24'h93895d,
24'h999b46,
24'h969a3c,
24'h5d5b10,
24'h4d4608,
24'h575316,
24'h928958,
24'h877960,
24'h390d22,
24'h6f0e69,
24'h7d017e,
24'h7d017e,
24'h7d017e,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f0081,
24'h7f0083,
24'h7e0082,
24'h7c007e,
24'h7d047f,
24'h6c175c,
24'h7c6746,
24'h849337,
24'hb3c762,
24'hbccd6a,
24'h8d9240,
24'h908f4d,
24'h909262,
24'h241904,
24'h360e19,
24'h340d0d,
24'h555316,
24'h8f9b42,
24'h848d37,
24'h8b9339,
24'hc7d270,
24'h979d41,
24'h827e38,
24'h524719,
24'h2b1504,
24'h927f67,
24'h8c8a46,
24'h93983e,
24'h8f933e,
24'h595b09,
24'h959348,
24'h908351,
24'h2f130f,
24'h4f1442,
24'h710b6e,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f0081,
24'h7f0083,
24'h7e0084,
24'h7e0082,
24'h7c0281,
24'h6c1364,
24'h93786a,
24'hc4cb86,
24'hb7c770,
24'hc1d173,
24'hced37a,
24'h8d8943,
24'h898261,
24'h290d16,
24'h5c1a52,
24'h602447,
24'h948d57,
24'hb8ca6e,
24'h869142,
24'h889140,
24'hbcc965,
24'h898e37,
24'h948757,
24'h5f4434,
24'h4c2931,
24'h270c0c,
24'h676437,
24'h89924e,
24'h6b702b,
24'h8d8d4b,
24'h746a30,
24'h9c8067,
24'h380524,
24'h5c0e5a,
24'h750776,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f0081,
24'h7f0083,
24'h7e0085,
24'h7e0084,
24'h7c0281,
24'h6c1169,
24'h532d3f,
24'h706b4a,
24'hc3ca8c,
24'h8c9844,
24'hc7cc6c,
24'h969147,
24'h837563,
24'h26001d,
24'h68145d,
24'h671e4c,
24'h867e4b,
24'hbcd172,
24'hb3c46f,
24'hbfd077,
24'hb8c861,
24'h909248,
24'h2e110f,
24'h56274d,
24'h5b2651,
24'h502c46,
24'hc4c7b9,
24'h334222,
24'hd4d6bd,
24'h493c2c,
24'heac9c5,
24'h612a47,
24'h600b5d,
24'h6a0273,
24'h79027c,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f0081,
24'h7f0083,
24'h820085,
24'h800085,
24'h7c0281,
24'h700d6f,
24'h5f2956,
24'hfff8fe,
24'h4d422b,
24'hffffe3,
24'h584f13,
24'h94825a,
24'h300a1c,
24'h5a1954,
24'h761569,
24'h6b194d,
24'h5d4b27,
24'hbbc67c,
24'h848f4e,
24'hbbc586,
24'h8e934e,
24'h968664,
24'h2f0022,
24'h5d1661,
24'h5e0f5e,
24'h541254,
24'h200323,
24'h18061b,
24'h250723,
24'h2f0025,
24'h3e002f,
24'h68145d,
24'h720879,
24'h7a0386,
24'h7b0081,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f0081,
24'h810083,
24'h880085,
24'h880084,
24'h80027f,
24'h760a72,
24'h61115e,
24'h360030,
24'h220019,
24'h2c0921,
24'h260215,
24'h370528,
24'h68175f,
24'h740f6a,
24'h770c64,
24'h78235c,
24'hfffaf5,
24'h4a4022,
24'hfffff3,
24'h453b31,
24'hfff3f5,
24'h370723,
24'h62155d,
24'h6e0a6e,
24'h760476,
24'h760476,
24'h6c0b6d,
24'h680d6a,
24'h6c0c6b,
24'h700a6d,
24'h74096e,
24'h760673,
24'h7a017b,
24'h7c0080,
24'h7d007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f0081,
24'h810083,
24'h880085,
24'h880084,
24'h80027f,
24'h780777,
24'h6f0e70,
24'h620f65,
24'h58105e,
24'h56145f,
24'h571161,
24'h600b66,
24'h7a0a78,
24'h810574,
24'h81096c,
24'h76115d,
24'h440029,
24'h35051f,
24'h2b0020,
24'h30002d,
24'h390036,
24'h651461,
24'h6e0b6d,
24'h780378,
24'h800080,
24'h820083,
24'h800080,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f0081,
24'h7f0081,
24'h800084,
24'h800084,
24'h7c0281,
24'h78047d,
24'h6f0374,
24'h700977,
24'h6e0e76,
24'h6e0a75,
24'h78097f,
24'h810882,
24'h82007b,
24'h88027c,
24'h820071,
24'h840774,
24'h7c0b6f,
24'h7b1172,
24'h760c6f,
24'h77096f,
24'h750570,
24'h780575,
24'h7a0378,
24'h7c017b,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7c007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7d0081,
24'h7c0084,
24'h7c0182,
24'h7c0182,
24'h7a0281,
24'h7f0785,
24'h77027e,
24'h75007b,
24'h79017f,
24'h78007c,
24'h850085,
24'h7f007a,
24'h890180,
24'h84007a,
24'h86007f,
24'h7e007b,
24'h7e007b,
24'h81007d,
24'h8a0686,
24'h7c007b,
24'h830280,
24'h7e007d,
24'h7e007d,
24'h7e007d,
24'h7c007d,
24'h7c007e,
24'h7c007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7e007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d0081,
24'h7c0182,
24'h7c0182,
24'h7c0182,
24'h7e0084,
24'h7e0084,
24'h800085,
24'h800085,
24'h800084,
24'h81007e,
24'h81017c,
24'h7f007f,
24'h7e0082,
24'h7c0080,
24'h7e0080,
24'h80007e,
24'h7e007d,
24'h79027c,
24'h77037c,
24'h79027c,
24'h79027e,
24'h7b017e,
24'h7d017e,
24'h7f007e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7d007f,
24'h7d007f,
24'h800082,
24'h800082,
24'h800082,
24'h800084,
24'h820084,
24'h820085,
24'h820085,
24'h820082,
24'h81027b,
24'h7f027b,
24'h7d017e,
24'h7d0081,
24'h7c0080,
24'h7c007e,
24'h7e007b,
24'h7c017b,
24'h77027e,
24'h75027f,
24'h75027f,
24'h77017f,
24'h7b007f,
24'h7d017e,
24'h7d017e,
24'h7f007e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f0081,
24'h810081,
24'h860082,
24'h880082,
24'h860082,
24'h840081,
24'h82017f,
24'h82017f,
24'h80027d,
24'h80027d,
24'h7d027c,
24'h7d017e,
24'h81007e,
24'h83007e,
24'h82007b,
24'h800179,
24'h7c0376,
24'h7a0279,
24'h790084,
24'h790089,
24'h790087,
24'h7b0084,
24'h7b0081,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f0081,
24'h810081,
24'h860082,
24'h880082,
24'h860081,
24'h84017f,
24'h82027d,
24'h80037c,
24'h80037c,
24'h7e047c,
24'h7d017e,
24'h7d007f,
24'h81007e,
24'h83007e,
24'h82007b,
24'h800178,
24'h7c0376,
24'h7c017b,
24'h7d0086,
24'h7d0089,
24'h7d0087,
24'h7d0086,
24'h7d0083,
24'h7d007f,
24'h7d017e,
24'h7d017e,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h820081,
24'h820081,
24'h820081,
24'h820081,
24'h80027f,
24'h80027f,
24'h80027f,
24'h80027f,
24'h800181,
24'h800181,
24'h800181,
24'h820081,
24'h81007e,
24'h7f007e,
24'h7f017c,
24'h7f007e,
24'h7f0081,
24'h7f0083,
24'h7f0083,
24'h7f0081,
24'h7f0081,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h800181,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
24'h7f007f,
};

    always_ff @(posedge clk) begin
        o_rd_data[0][2] <= bulbasaur_rom_buf[i_rd_addr][3*bpp_p-1-:8];
        o_rd_data[0][1] <= bulbasaur_rom_buf[i_rd_addr][2*bpp_p-1-:8];
        o_rd_data[0][0] <= bulbasaur_rom_buf[i_rd_addr][1*bpp_p-1-:8];

        o_rd_data[1][2] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][3*bpp_p-1-:8];
        o_rd_data[1][1] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][2*bpp_p-1-:8];
        o_rd_data[1][0] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][1*bpp_p-1-:8];
    end
endmodule