module bulbasaur_rom #(
    parameter hpixel_p = 64,
    parameter vpixel_p = 64,
    parameter bpp_p = 8,
    parameter segments_p = 2,
    localparam frame_size_p = hpixel_p*vpixel_p,
    localparam addr_width_p = $clog2(frame_size_p)
    ) (

    // Clock and reset
    input logic clk,
    input logic rst_n,

    /* Pixel read interface */
    input logic [addr_width_p-1:0] i_rd_addr,
    output logic [segments_p-1:0][2:0][bpp_p-1:0] o_rd_data
    );

	localparam [frame_size_p-1:0][3*bpp_p-1:0] bulbasaur_rom_buf = {
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x80007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x80007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x80007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x80007f,
		0x81007f,
		0x82007f,
		0x83007f,
		0x82007f,
		0x7f007f,
		0x7d017f,
		0x7d017f,
		0x7e0080,
		0x7f0082,
		0x810081,
		0x810180,
		0x810180,
		0x800180,
		0x7f0280,
		0x7f0280,
		0x7f0280,
		0x800181,
		0x810082,
		0x810082,
		0x810082,
		0x810081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e017e,
		0x7e017d,
		0x7e007d,
		0x81007d,
		0x85007d,
		0x87007d,
		0x88007d,
		0x88007d,
		0x81007c,
		0x78027c,
		0x76027e,
		0x790081,
		0x7d0083,
		0x7e0082,
		0x7e007f,
		0x7f007d,
		0x7d027d,
		0x7c047f,
		0x7c0380,
		0x7c0381,
		0x7e0283,
		0x800185,
		0x810087,
		0x820088,
		0x820085,
		0x810080,
		0x81007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e017e,
		0x7e017d,
		0x7e007d,
		0x80007c,
		0x83007b,
		0x86007a,
		0x89007a,
		0x880079,
		0x7e0179,
		0x77037b,
		0x77027e,
		0x7a0081,
		0x7c0083,
		0x7e0082,
		0x7e007f,
		0x7d017d,
		0x7c027e,
		0x7d0280,
		0x7d0281,
		0x7e0182,
		0x800182,
		0x810085,
		0x820087,
		0x820088,
		0x820085,
		0x810080,
		0x81007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e017e,
		0x7e017d,
		0x7f007c,
		0x7f0079,
		0x800276,
		0x800275,
		0x800276,
		0x7c027a,
		0x7a007d,
		0x7b007d,
		0x7e007c,
		0x80007d,
		0x80007d,
		0x7d017e,
		0x7a0280,
		0x7d0182,
		0x830082,
		0x840082,
		0x840082,
		0x840081,
		0x830081,
		0x820081,
		0x820081,
		0x810080,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e017e,
		0x7e017c,
		0x7e0279,
		0x7d0278,
		0x7c0377,
		0x7c0377,
		0x7c017c,
		0x7d007f,
		0x7f007f,
		0x80007c,
		0x81007c,
		0x81007d,
		0x7e0080,
		0x7b0181,
		0x800082,
		0x850081,
		0x860081,
		0x850080,
		0x84007e,
		0x83007d,
		0x82017c,
		0x82017c,
		0x82017c,
		0x81007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007d,
		0x7e007c,
		0x7d007c,
		0x7d007d,
		0x7d007e,
		0x7d007e,
		0x7f0181,
		0x7e017e,
		0x810483,
		0x820385,
		0x7c007f,
		0x7c007d,
		0x7e0082,
		0x7e0084,
		0x7e0086,
		0x7e0184,
		0x7e0081,
		0x810081,
		0x7e0079,
		0x7f007a,
		0x7d0077,
		0x81037b,
		0x85057f,
		0x81017a,
		0x82017c,
		0x83017c,
		0x84007c,
		0x80007d,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007c,
		0x7e007d,
		0x7e007d,
		0x7e007e,
		0x7c007d,
		0x7a017c,
		0x78037b,
		0x76047a,
		0x76077d,
		0x770a7d,
		0x780e7e,
		0x770e7f,
		0x760883,
		0x740284,
		0x770086,
		0x7c0186,
		0x7f0283,
		0x840781,
		0x7d0776,
		0x780a70,
		0x790b71,
		0x780672,
		0x780373,
		0x80047a,
		0x82017c,
		0x84007f,
		0x83007f,
		0x81007f,
		0x81007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007e,
		0x7e007e,
		0x7f007e,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x800080,
		0x820082,
		0x820081,
		0x7d007d,
		0x740574,
		0x6e1170,
		0x49004c,
		0x330036,
		0x2a0030,
		0x240033,
		0x27003e,
		0x41005b,
		0x6a0d80,
		0x710583,
		0x790581,
		0x760875,
		0x6d0d64,
		0x69125e,
		0x66135d,
		0x681062,
		0x6e0e6a,
		0x740a72,
		0x7a057b,
		0x810182,
		0x850088,
		0x850086,
		0x830080,
		0x81007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007c,
		0x7d007c,
		0x780379,
		0x75077a,
		0x750978,
		0x740975,
		0x730b72,
		0x740a73,
		0x790479,
		0x7b027b,
		0x750575,
		0x6c116e,
		0x34003f,
		0x9980a2,
		0x797283,
		0x878691,
		0x75818d,
		0x76818e,
		0xad8ebe,
		0x570a71,
		0x6a0979,
		0x6f1177,
		0x520d59,
		0x26002f,
		0x1f0027,
		0x1f0025,
		0x240029,
		0x3c0040,
		0x6b106d,
		0x77077b,
		0x810183,
		0x85008a,
		0x850087,
		0x830080,
		0x81007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x80007b,
		0x86027c,
		0x800577,
		0x6b1070,
		0x3c0048,
		0x31003a,
		0x29002b,
		0x280225,
		0x24001f,
		0x490647,
		0x620c63,
		0x691165,
		0x410343,
		0x423d60,
		0x68939b,
		0x76ada7,
		0x74a9a0,
		0x6faea4,
		0x5e9494,
		0x4e4473,
		0x5b1273,
		0x681671,
		0x410c4a,
		0x352e52,
		0x315569,
		0x51737e,
		0x94a1ab,
		0x565a69,
		0xc6abc6,
		0x55115b,
		0x760875,
		0x83017f,
		0x850083,
		0x850083,
		0x83007f,
		0x81007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7e017b,
		0x7b0072,
		0x6d0769,
		0x481258,
		0x9f8ebc,
		0x44455e,
		0x879198,
		0x40534b,
		0x77837d,
		0x6d5873,
		0x4e1e55,
		0x59235c,
		0x230631,
		0x305463,
		0x56afa6,
		0x70cdbd,
		0x74c7b6,
		0x71cbb7,
		0x5ba89f,
		0x40416c,
		0x59146c,
		0x48084e,
		0x362544,
		0x527683,
		0x50a2a5,
		0x5db5ae,
		0x6fb1a9,
		0x7ba6a5,
		0x606978,
		0x481a54,
		0x730b73,
		0x83007e,
		0x84007e,
		0x85007f,
		0x83007f,
		0x81007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x80007e,
		0x7b0479,
		0x680a66,
		0x380142,
		0x55537c,
		0x5a8194,
		0x4b8086,
		0x4d8885,
		0x478479,
		0x578681,
		0x283042,
		0x2a193f,
		0x3c3459,
		0x445a71,
		0x3d7f83,
		0x52b5a9,
		0x59b6aa,
		0x4a998e,
		0x62bbaa,
		0x6ab9b0,
		0x51597c,
		0x541963,
		0x390b42,
		0x34384c,
		0x59898f,
		0x58aaab,
		0x78d6cd,
		0x6ac4b4,
		0x7cc8bc,
		0x729fa5,
		0x604b7b,
		0x6d086e,
		0x83007e,
		0x83007e,
		0x84007e,
		0x83007f,
		0x81007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x80007e,
		0x760776,
		0x55135c,
		0x13022a,
		0x46677c,
		0x4c8f95,
		0x217170,
		0x2e807c,
		0x419891,
		0x3f8787,
		0x4f6f7d,
		0x252f48,
		0x132e41,
		0x346c76,
		0x3f908f,
		0x5dbfb5,
		0x52aea4,
		0x33867e,
		0x459d91,
		0x3d8c84,
		0x1c344d,
		0x1d0337,
		0x110327,
		0x2c474e,
		0x669d9d,
		0x4c9696,
		0x5ab4ab,
		0x6ed2be,
		0x5cbdaa,
		0x4b9490,
		0x53517b,
		0x680a6e,
		0x82017e,
		0x80007d,
		0x83007d,
		0x83007f,
		0x81007f,
		0x7f007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7e017d,
		0x7e017d,
		0x7f007e,
		0x720b75,
		0x350a45,
		0x424a61,
		0x57838e,
		0x337176,
		0x0a4d52,
		0x135e5f,
		0x338e8b,
		0x439c99,
		0x63979f,
		0x223d4d,
		0x08313c,
		0x327377,
		0x3b8c8b,
		0x5dbcb6,
		0x68cfc6,
		0x3ea69c,
		0x3d9b92,
		0x24716c,
		0x164f56,
		0x3d6775,
		0x3c696e,
		0x26574f,
		0x134742,
		0x256d6c,
		0x52a89e,
		0x6fd5c0,
		0x52bba5,
		0x2d827a,
		0x404c71,
		0x5f0c6c,
		0x7e037e,
		0x7e027c,
		0x880684,
		0x81007d,
		0x80007e,
		0x7e007e,
		0x7d007e,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7e017d,
		0x7e017d,
		0x80007e,
		0x710d77,
		0x1a0132,
		0x4d6676,
		0x5f8e96,
		0x225b61,
		0x0d444c,
		0x0b4b50,
		0x247c7a,
		0x3b9b96,
		0x569c9f,
		0x1a363e,
		0x002c30,
		0x347b7b,
		0x419291,
		0x3e9c98,
		0x59c3be,
		0x68d8d1,
		0x32908a,
		0x1c6664,
		0x3d8b85,
		0x489e90,
		0x54a190,
		0x4c8d7d,
		0x427d74,
		0x327270,
		0x2a7a71,
		0x60c2af,
		0x6cd5bf,
		0x65bcb1,
		0x7f91b3,
		0x7e3793,
		0x740379,
		0x790077,
		0x870382,
		0x82007e,
		0x80007e,
		0x7d007e,
		0x7d007e,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7e017d,
		0x7e017d,
		0x80007e,
		0x700c78,
		0x1d053d,
		0x4f6e83,
		0x548893,
		0x1a575e,
		0x114d52,
		0x0c4d50,
		0x2c817c,
		0x3d9d93,
		0x1e5e58,
		0x2a5856,
		0x397976,
		0x1c6a66,
		0x257e7b,
		0x359392,
		0x3e989b,
		0x53a9ae,
		0x459497,
		0x46908e,
		0x306c5f,
		0x093720,
		0x0d3f28,
		0x103c2c,
		0x14413a,
		0x073736,
		0x002b24,
		0x0f4633,
		0x185641,
		0x366c65,
		0x7c8caf,
		0x692b85,
		0x6d0378,
		0x7d017b,
		0x7e0077,
		0x83007f,
		0x80007e,
		0x7d007f,
		0x7d007e,
		0x7f007f,
		0x7f007e,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7e017d,
		0x7e017d,
		0x80007e,
		0x700c78,
		0x210141,
		0x576e8b,
		0x528796,
		0x387b82,
		0x115356,
		0x276c6b,
		0x3e9087,
		0x439d8f,
		0x0e574b,
		0x2e7269,
		0x47958f,
		0x1e746c,
		0x1f7a75,
		0x3a9294,
		0x4a98a1,
		0x2a606e,
		0x123841,
		0x153f41,
		0x275148,
		0x4b6754,
		0x4f6251,
		0x565e55,
		0x535859,
		0x4f555e,
		0x4e585c,
		0x495f59,
		0x496960,
		0x355655,
		0x151936,
		0x2d0550,
		0x641478,
		0x760977,
		0x7e0378,
		0x82007d,
		0x80007f,
		0x7d0080,
		0x7c0080,
		0x80007e,
		0x80007d,
		0x800080,
		0x800080,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e007e,
		0x7e017d,
		0x7e017d,
		0x7f007e,
		0x730977,
		0x3f0d51,
		0x3d3f63,
		0x4e798a,
		0x4e9297,
		0x37807d,
		0x458f89,
		0x4b9a8f,
		0x36887b,
		0x2d7c70,
		0x39877d,
		0x3e958b,
		0x338e85,
		0x408f8e,
		0x27636b,
		0x133842,
		0x275762,
		0x336c78,
		0x2e606b,
		0x56757a,
		0x807d7d,
		0x9e787a,
		0xc7848c,
		0xcf7b8c,
		0xd27d96,
		0xc3708c,
		0x914962,
		0x724559,
		0x6e6370,
		0x4f5166,
		0x414267,
		0x1b053a,
		0x43054c,
		0x781675,
		0x7e0075,
		0x83007e,
		0x77007c,
		0x75007b,
		0x80007d,
		0x82007e,
		0x830084,
		0x830085,
		0x800080,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e017d,
		0x7e017d,
		0x7f017e,
		0x750777,
		0x5d1465,
		0x432759,
		0x597387,
		0x549294,
		0x4b938f,
		0x28746d,
		0x1d675e,
		0x358076,
		0x4e9990,
		0x44948c,
		0x3d968e,
		0x429c95,
		0x2c7374,
		0x2b5e67,
		0x38646c,
		0x427f86,
		0x4d97a2,
		0x40828f,
		0x45626d,
		0x5b474f,
		0x7f3d47,
		0xa13b4a,
		0xa9334a,
		0xa72e4c,
		0xa02348,
		0x8b143b,
		0x60112e,
		0x4c3140,
		0x4e565e,
		0x5e757e,
		0x4a596d,
		0x4f3e63,
		0x571c5e,
		0x73096f,
		0x81067e,
		0x7b0481,
		0x75007a,
		0x80007c,
		0x83007f,
		0x840088,
		0x840089,
		0x810082,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e017d,
		0x7e017d,
		0x7e017d,
		0x79057a,
		0x68066f,
		0x5a1d6a,
		0x474a65,
		0x50817d,
		0x559791,
		0x1b5f5c,
		0x0b4a46,
		0x23615b,
		0x448b86,
		0x499a93,
		0x419690,
		0x277a77,
		0x236d6d,
		0x46878a,
		0x5c9b9f,
		0x58999c,
		0x3b8283,
		0x71b0b4,
		0x608182,
		0x0b0906,
		0x1b0e09,
		0x361817,
		0x523235,
		0x71545a,
		0x987b85,
		0x9d838f,
		0x828184,
		0x708c87,
		0x5c7373,
		0x33323f,
		0x6f707e,
		0xc7d2dd,
		0x5a4d78,
		0x4e1361,
		0x650770,
		0x7d0983,
		0x7c017f,
		0x7c027c,
		0x7f0080,
		0x820088,
		0x840087,
		0x810081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e017d,
		0x7e017d,
		0x7e017d,
		0x7c037c,
		0x6d0073,
		0x651c71,
		0x1f1b30,
		0x1d4b3a,
		0x498a7f,
		0x448584,
		0x1d5858,
		0x0a4443,
		0x307573,
		0x449490,
		0x459593,
		0x247271,
		0x2d7c7a,
		0x4d9b9a,
		0x316668,
		0x1a3d3f,
		0x0d453e,
		0x417e72,
		0x719d8f,
		0x5c7a6a,
		0x4f7866,
		0x548775,
		0x609e8c,
		0x72bca8,
		0x68b5a2,
		0x5daa97,
		0x88ddc7,
		0x73c8b1,
		0x6d9b93,
		0x837e8b,
		0x817b88,
		0x5f7478,
		0x2b3a52,
		0x65578b,
		0x4e1368,
		0x74077b,
		0x7e017d,
		0x7b037d,
		0x7a0280,
		0x7f0086,
		0x810085,
		0x800081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7d017d,
		0x800480,
		0x7e027f,
		0x740173,
		0x721671,
		0x3a093d,
		0x34453a,
		0x2f6e43,
		0x1d6951,
		0x45918d,
		0x44898e,
		0x307379,
		0x408588,
		0x4a9494,
		0x449693,
		0x358c88,
		0x388c88,
		0x2b7777,
		0x285e63,
		0x2e5054,
		0x436a61,
		0x628773,
		0x90ac9a,
		0xb3cfc3,
		0x98cabb,
		0x80d2be,
		0x72d7bf,
		0x6ad9bf,
		0x4fc0a6,
		0x48b89e,
		0x68dbbf,
		0x5cccb0,
		0x65bca7,
		0x9dd3c8,
		0x99b5b4,
		0x6c757b,
		0x596271,
		0x263150,
		0x47276a,
		0x720a7a,
		0x80017f,
		0x7a027e,
		0x79037f,
		0x7d0184,
		0x7e0084,
		0x7f0081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f0481,
		0x800581,
		0x800481,
		0x770d77,
		0x4e104a,
		0x3d313a,
		0x538054,
		0x51a162,
		0x2e835d,
		0x1e7164,
		0x1e6e6d,
		0x3f8c90,
		0x4e9699,
		0x4b9092,
		0x409491,
		0x399891,
		0x3f9893,
		0x368281,
		0x417e83,
		0x79a1a9,
		0xa0adaa,
		0xada296,
		0x947d79,
		0x675d5f,
		0x618581,
		0x68bdad,
		0x66d4bc,
		0x5bd1b6,
		0x5bd2b9,
		0x64d6bf,
		0x5dd3b9,
		0x5bd4b7,
		0x60d8b8,
		0x61ccad,
		0x5e9283,
		0x6c5c62,
		0x786d7a,
		0x4c6473,
		0x514275,
		0x721079,
		0x7f007c,
		0x7a027f,
		0x7a037f,
		0x7b0282,
		0x7d0082,
		0x7e0080,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7d017e,
		0x7d017e,
		0x7e007f,
		0x7e007f,
		0x7f0480,
		0x80057f,
		0x820482,
		0x761377,
		0x1f001d,
		0x496248,
		0x519055,
		0x489858,
		0x348254,
		0x257053,
		0x24745c,
		0x1a6c5b,
		0x3a857e,
		0x4c9394,
		0x3a8989,
		0x39948d,
		0x38988f,
		0x3c9692,
		0x67a7ac,
		0xc1d9e2,
		0xd9b7c3,
		0xd17e8c,
		0xce8fa2,
		0x7b576d,
		0x43434e,
		0x62a89e,
		0x70d8bf,
		0x70e2c1,
		0x77e5ca,
		0x7de3d1,
		0x78e2cf,
		0x6ee3c7,
		0x6be3c1,
		0x5cc2a2,
		0x61897d,
		0x90707f,
		0x674553,
		0xcce0e5,
		0x534871,
		0x67086e,
		0x7c007c,
		0x7d017f,
		0x7c017f,
		0x7b0280,
		0x7b0280,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7c027d,
		0x7d027d,
		0x7e0080,
		0x7e0080,
		0x7a017b,
		0x820a82,
		0x7d047c,
		0x540653,
		0x393539,
		0x487f4a,
		0x489150,
		0x2e7a3d,
		0x347c47,
		0x418958,
		0x469766,
		0x257c50,
		0x1b6a51,
		0x3f8881,
		0x2b7470,
		0x2f807a,
		0x3c9d93,
		0x2d918a,
		0x7dc1c6,
		0xf0ffff,
		0xd495aa,
		0xa82744,
		0xf19ac2,
		0xd0a3c8,
		0x604559,
		0x6fa9a2,
		0x89e8ce,
		0x8bf4d1,
		0x7fe1c7,
		0x61b6ac,
		0x6ecdbe,
		0x88f7dc,
		0x83f0cf,
		0x6ec2a6,
		0x88a29b,
		0xf8d6eb,
		0x89556a,
		0xdddfeb,
		0x59436f,
		0x65036a,
		0x7d007c,
		0x7e007f,
		0x7c017f,
		0x7b027f,
		0x7b027f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x800180,
		0x800180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e017e,
		0x7b017b,
		0x7d007c,
		0x810082,
		0x820084,
		0x7a007b,
		0x7c097b,
		0x720c6f,
		0x34002f,
		0x526750,
		0x4f974f,
		0x46924b,
		0x236d2e,
		0x408f52,
		0x3d9254,
		0x358f4d,
		0x3c9655,
		0x2b7e4d,
		0x276f54,
		0x0e4839,
		0x286860,
		0x439892,
		0x3d9793,
		0x468a8f,
		0xbbd2d5,
		0xe1c2cc,
		0x9b3657,
		0xaa3c69,
		0xb07095,
		0x847584,
		0x86c8bb,
		0x83e6c9,
		0x79ddbd,
		0x48a48e,
		0x308479,
		0x4eab9b,
		0x8bf6d8,
		0x82eac8,
		0x7ccfb2,
		0x98b4ab,
		0xbc98ac,
		0x864e72,
		0x88699a,
		0x612a74,
		0x700572,
		0x7d0078,
		0x7d027d,
		0x7c027e,
		0x7c027e,
		0x7d017e,
		0x7f007e,
		0x7f007e,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e017d,
		0x7b017a,
		0x7c007b,
		0x820083,
		0x840086,
		0x7c007e,
		0x730573,
		0x6a1464,
		0x2a0322,
		0x496c45,
		0x469544,
		0x358138,
		0x388043,
		0x378e4e,
		0x31924d,
		0x399a4c,
		0x399344,
		0x479956,
		0x236c3b,
		0x00270c,
		0x2e5c51,
		0x428b85,
		0x429490,
		0x135b5b,
		0x759a9d,
		0xffffff,
		0xbe85a4,
		0x6d1739,
		0x703f57,
		0x829496,
		0x91e3cf,
		0x6fd6b9,
		0x62c5ab,
		0x27826f,
		0x449a8e,
		0x71cdba,
		0x89efcf,
		0x81e6c1,
		0x80d8b6,
		0x9dc8b9,
		0x72616f,
		0x6c406e,
		0x4d1365,
		0x630c76,
		0x7b0379,
		0x80007a,
		0x7b037d,
		0x7a037d,
		0x7c027d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e017d,
		0x7b017a,
		0x7c007b,
		0x820083,
		0x840086,
		0x7b007e,
		0x740573,
		0x6a1365,
		0x2c0224,
		0x466947,
		0x47984d,
		0x23702c,
		0x3f8a4e,
		0x368d4f,
		0x36954f,
		0x3c9748,
		0x4fa151,
		0x5ead65,
		0x539e63,
		0x0a3613,
		0x305a4a,
		0x499588,
		0x339386,
		0x389287,
		0x498a86,
		0xacc6c8,
		0xc4bdc7,
		0x6b656e,
		0x5f7374,
		0x7db9ac,
		0x7bdcc3,
		0x76e3c5,
		0x72dabf,
		0x5cbaa6,
		0x7dd1c5,
		0x96edd9,
		0x8ae6c8,
		0x86e7c2,
		0x78dab4,
		0x80cab2,
		0x769697,
		0x4e3f69,
		0x672883,
		0x6a0579,
		0x80037d,
		0x7f0079,
		0x7b037c,
		0x7a037c,
		0x7c027d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007e,
		0x7c017b,
		0x7d007d,
		0x820083,
		0x840084,
		0x7c007d,
		0x770575,
		0x700f6b,
		0x30002d,
		0x526b59,
		0x4e9a5d,
		0x257537,
		0x37854a,
		0x3c8f51,
		0x419653,
		0x53a057,
		0x72b970,
		0x76c37a,
		0x77c485,
		0x5d926b,
		0x355c47,
		0x337f6b,
		0x42b19b,
		0x63d1bb,
		0x4aa794,
		0x4d9386,
		0x88c0b4,
		0x6db2a2,
		0x6fc7b0,
		0x8bf0d4,
		0x77e2c4,
		0x86f3d5,
		0x7ae5c9,
		0x63c4af,
		0x6dc3b4,
		0x74c8b4,
		0x8de3c5,
		0x8cebc6,
		0x7de9c1,
		0x79e0bf,
		0x7bc6bb,
		0x344364,
		0x652782,
		0x71057a,
		0x7f027b,
		0x7c0076,
		0x7c027b,
		0x7b037b,
		0x7c027d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x80007f,
		0x810180,
		0x810180,
		0x80007f,
		0x80007f,
		0x80007f,
		0x800080,
		0x7f017e,
		0x7f007f,
		0x830083,
		0x830083,
		0x7f007f,
		0x7a0379,
		0x760a73,
		0x4b0a4a,
		0x3d4346,
		0x48835a,
		0x226e3a,
		0x34844b,
		0x3e9151,
		0x53a360,
		0x7ac07b,
		0x80c47d,
		0x76c279,
		0x76c580,
		0xace6b8,
		0x406045,
		0x11533c,
		0x58c6ac,
		0x65d9bd,
		0x69d7ba,
		0x5dbfa4,
		0x45a188,
		0x59c4a6,
		0x76efcd,
		0x84f7d7,
		0x8bf1d5,
		0x79dcc1,
		0x4fb198,
		0x2f927c,
		0x2a8d79,
		0x4eab94,
		0x93eacb,
		0x8feec9,
		0x7febc3,
		0x82f0cd,
		0x75cdbf,
		0x3e5273,
		0x530e6a,
		0x79057d,
		0x7e007a,
		0x80007a,
		0x7d027b,
		0x7b037b,
		0x7d027d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x80007f,
		0x800080,
		0x830083,
		0x830083,
		0x820182,
		0x7f017e,
		0x7c047a,
		0x6d156d,
		0x14001d,
		0x456857,
		0x397b54,
		0x2b7d45,
		0x378949,
		0x63b36e,
		0x7dc581,
		0x7bc17b,
		0x7ece82,
		0x8cde94,
		0xa7e5b0,
		0x345738,
		0x18543b,
		0x5cbba2,
		0x66d3b5,
		0x65d8b4,
		0x6ad8b7,
		0x67d1b4,
		0x5dd6b4,
		0x66ebc5,
		0x81f7d6,
		0x7edec5,
		0x51a891,
		0x348d76,
		0x369983,
		0x33a38b,
		0x69d2b6,
		0x8fedcb,
		0x88e9c4,
		0x81e9c2,
		0x77dfbf,
		0x4fa397,
		0x536185,
		0x5e0d6e,
		0x7d027c,
		0x7f017b,
		0x80007b,
		0x7f017b,
		0x7d027b,
		0x7e017d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810181,
		0x810181,
		0x820181,
		0x820082,
		0x820082,
		0x820082,
		0x820082,
		0x820182,
		0x820181,
		0x740a75,
		0x390c40,
		0x354045,
		0x538a6e,
		0x20713d,
		0x2a7e3d,
		0x5db069,
		0x75c37f,
		0x73c17a,
		0x86db8a,
		0x94e898,
		0x9bdda3,
		0x64926e,
		0x2d5c44,
		0x5a9a85,
		0x74cbb0,
		0x6fd9b5,
		0x72debc,
		0x73dec0,
		0x65ddbc,
		0x5bdeb9,
		0x7af2d0,
		0x63caad,
		0x2e8c73,
		0x37937b,
		0x40a38c,
		0x65d0b9,
		0x8cf1d6,
		0x90efcc,
		0x8ef1ca,
		0x7ce7be,
		0x56bd9c,
		0x47968b,
		0x666d92,
		0x64096e,
		0x81007d,
		0x7f007c,
		0x7f007c,
		0x7f007c,
		0x7f017c,
		0x7e017d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x820082,
		0x820082,
		0x820082,
		0x820082,
		0x820082,
		0x820082,
		0x820082,
		0x830083,
		0x860086,
		0x7b037c,
		0x651c67,
		0x1a0724,
		0x4f7264,
		0x377d51,
		0x257537,
		0x5aae67,
		0x6dc47e,
		0x68c078,
		0x80d987,
		0x90e593,
		0x8fd798,
		0xb1ebc1,
		0x3c6048,
		0x4a6e5e,
		0x94d6bd,
		0x8ae6c2,
		0x96f7d6,
		0x6ccbaf,
		0x50bb9d,
		0x63d9b7,
		0x71e3c3,
		0x71dbbe,
		0x59b9a0,
		0x5cb4a0,
		0x72c7b9,
		0x9bede2,
		0x87d5c6,
		0x6bb9a0,
		0x76ceb0,
		0x7ae0bd,
		0x60c0a6,
		0x94dad5,
		0x63608a,
		0x680770,
		0x83007e,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7f007d,
		0x7e017d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x820081,
		0x820081,
		0x820081,
		0x820081,
		0x820081,
		0x820081,
		0x820082,
		0x830083,
		0x850085,
		0x80017f,
		0x750f73,
		0x420444,
		0x413d4f,
		0x59806d,
		0x347042,
		0x5da86a,
		0x68c17d,
		0x63c17a,
		0x7cd68b,
		0x8bdd93,
		0x90da9c,
		0xa2e3b3,
		0x325e3d,
		0x4f7962,
		0xaeefd3,
		0x80d1af,
		0x5fb496,
		0x287d63,
		0x1f775c,
		0x57b397,
		0x57ad95,
		0x6cb7a7,
		0x87bebd,
		0x8db2bf,
		0x91aec1,
		0x95aec3,
		0x73889d,
		0x2c4453,
		0x436e75,
		0x84c5c5,
		0xa9ecef,
		0xa1d0e1,
		0x6a5b92,
		0x690571,
		0x82007e,
		0x7f007d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7e017e,
		0x7e017e,
		0x7f007e,
		0x7f007e,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x820082,
		0x820082,
		0x810081,
		0x820180,
		0x7f007a,
		0x760e73,
		0x3a073f,
		0x45434f,
		0x3b5a43,
		0x599363,
		0x66b778,
		0x62c07b,
		0x79d18a,
		0x92df9e,
		0x7ec88c,
		0x74bd86,
		0x316e3f,
		0x326941,
		0x67a884,
		0x4a9472,
		0x287353,
		0x38856a,
		0x4a9177,
		0x548f7a,
		0x5b867d,
		0x485d67,
		0x484163,
		0x56336b,
		0x5e3271,
		0x633577,
		0x5f2f71,
		0x4f2363,
		0x3c2861,
		0x444f7d,
		0x90a6d0,
		0x808bbb,
		0x64408b,
		0x6d0576,
		0x80007e,
		0x7e017d,
		0x7e017d,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x820081,
		0x820081,
		0x810180,
		0x810080,
		0x880389,
		0x7e0782,
		0x681b6c,
		0x1f0024,
		0x303c35,
		0x4b7852,
		0x68ac73,
		0x71c17e,
		0x64b46b,
		0x73be76,
		0x68b36c,
		0x57a25f,
		0x5da96c,
		0x3b7a42,
		0x225e2b,
		0x6ab283,
		0xa4eebd,
		0x9ee5b8,
		0xa6ddbd,
		0xabcbbf,
		0x8b8b9a,
		0x603c68,
		0x57185d,
		0x5d0961,
		0x650a6a,
		0x670b6d,
		0x6b0f70,
		0x691071,
		0x5f1974,
		0x4a1f70,
		0x3d1c69,
		0x401667,
		0x571171,
		0x76067c,
		0x80007e,
		0x7e017e,
		0x7e017e,
		0x7f007e,
		0x7f007e,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x810180,
		0x800083,
		0x80028b,
		0x770282,
		0x6b0f70,
		0x2e0030,
		0x444248,
		0x4b6f52,
		0x72aa75,
		0x7cbc7a,
		0x61a458,
		0x4c9040,
		0x81c679,
		0xa3e79f,
		0xa0e4a0,
		0xa2e6a8,
		0xa2e5ac,
		0xa0e1aa,
		0x9edea3,
		0x99d099,
		0x9dc0a1,
		0x888b90,
		0x5c2f5d,
		0x63095b,
		0x7c0d74,
		0x810d7e,
		0x800b81,
		0x7c097d,
		0x790679,
		0x7a057b,
		0x720678,
		0x6c0d7b,
		0x620975,
		0x721283,
		0x790d81,
		0x7b017e,
		0x80007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x800180,
		0x7f0180,
		0x82068a,
		0x75007c,
		0x751176,
		0x40013e,
		0x635667,
		0x48644d,
		0x609461,
		0x558f4d,
		0x77aa6d,
		0x7fa774,
		0x6f9566,
		0x83aa7e,
		0x8aaf8a,
		0x8bae90,
		0x93b79c,
		0x97baa3,
		0x9db9a2,
		0x7c8779,
		0x625061,
		0x653267,
		0x630e64,
		0x780676,
		0x840580,
		0x860583,
		0x830484,
		0x7a017e,
		0x77017c,
		0x7e0281,
		0x79007d,
		0x7b0180,
		0x78017e,
		0x810684,
		0x79007b,
		0x7f0080,
		0x7f0080,
		0x7f0080,
		0x7f0080,
		0x7f0080,
		0x7f0080,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7d027c,
		0x780375,
		0x73086b,
		0x580851,
		0x5d3d5e,
		0x36463d,
		0x507d52,
		0x50824c,
		0x738c6f,
		0x5b5c59,
		0x40393f,
		0x423c44,
		0x3f3846,
		0x50485c,
		0x655c75,
		0x695d7c,
		0x6d507b,
		0x622c6a,
		0x5c0960,
		0x730773,
		0x7b0782,
		0x790284,
		0x7d0083,
		0x7f0082,
		0x7e0083,
		0x7c0185,
		0x7b0286,
		0x790284,
		0x7b0082,
		0x820083,
		0x810084,
		0x7f0081,
		0x7f0082,
		0x7f0081,
		0x7f0081,
		0x7f0081,
		0x7f0081,
		0x7e0081,
		0x7e0081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e017e,
		0x7d027a,
		0x7a0478,
		0x780776,
		0x6e0d6c,
		0x410041,
		0x1c001d,
		0x6f6a6d,
		0x5b6055,
		0x4d3748,
		0x52224e,
		0x551f52,
		0x501a51,
		0x511a57,
		0x50195b,
		0x4a1259,
		0x541564,
		0x62116e,
		0x6b0571,
		0x770379,
		0x800380,
		0x800284,
		0x7e0185,
		0x7f0086,
		0x830086,
		0x830085,
		0x800084,
		0x7c0184,
		0x790383,
		0x7d0082,
		0x850082,
		0x830082,
		0x7d0081,
		0x7d0081,
		0x7f0081,
		0x7f0081,
		0x7f0081,
		0x7f0081,
		0x7e0081,
		0x7e0081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7c027e,
		0x7b037e,
		0x790381,
		0x780381,
		0x710070,
		0x710969,
		0x6b2062,
		0x602356,
		0x621356,
		0x700f65,
		0x79136f,
		0x710b6a,
		0x730d72,
		0x710974,
		0x68006f,
		0x710479,
		0x7e0381,
		0x850085,
		0x7f017e,
		0x750173,
		0x790177,
		0x7f007d,
		0x840083,
		0x850088,
		0x870086,
		0x860080,
		0x81017e,
		0x7a027e,
		0x7e017e,
		0x85007e,
		0x82007e,
		0x79037e,
		0x79027f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7c017f,
		0x7b0280,
		0x7c0184,
		0x7e0086,
		0x80007e,
		0x810077,
		0x74036b,
		0x730e6b,
		0x76076c,
		0x7d0472,
		0x7e0275,
		0x7a0074,
		0x7c0078,
		0x7e017d,
		0x800283,
		0x850689,
		0x8a038a,
		0x8b0088,
		0x80007f,
		0x7c047b,
		0x81057e,
		0x80007c,
		0x830081,
		0x840085,
		0x860084,
		0x86007f,
		0x81017d,
		0x7c027d,
		0x7e017d,
		0x83007d,
		0x80017d,
		0x79047d,
		0x79037f,
		0x7d017f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7c017f,
		0x7c017f,
		0x7e0080,
		0x7f0080,
		0x810080,
		0x80007d,
		0x7d027b,
		0x7b0378,
		0x7c027a,
		0x7d007c,
		0x7e017c,
		0x7f017d,
		0x7e017e,
		0x7e007e,
		0x7e007f,
		0x7e007f,
		0x800080,
		0x820181,
		0x800180,
		0x7e007e,
		0x7e007d,
		0x80007e,
		0x800080,
		0x800080,
		0x81007f,
		0x82007f,
		0x80007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7d017f,
		0x7d017f,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f0080,
		0x7f0080,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e0081,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7c017f,
		0x7c017f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7c017f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7e007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007d,
		0x7f007d,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007d,
		0x81007d,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x7f007f,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007d,
		0x81007f,
		0x81007f,
		0x81007f,
		0x81007f,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081,
		0x810081
	};

    always_ff @(posedge clk) begin
        o_rd_data[0][2] <= bulbasaur_rom_buf[i_rd_addr][3*bpp_p-1-:8];
        o_rd_data[0][1] <= bulbasaur_rom_buf[i_rd_addr][2*bpp_p-1-:8];
        o_rd_data[0][0] <= bulbasaur_rom_buf[i_rd_addr][1*bpp_p-1-:8];

        o_rd_data[1][2] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][3*bpp_p-1-:8];
        o_rd_data[1][1] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][2*bpp_p-1-:8];
        o_rd_data[1][0] <= bulbasaur_rom_buf[i_rd_addr+frame_size_p/2][1*bpp_p-1-:8];
    end
endmodule